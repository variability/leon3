------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2006, Gaisler Research AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING. 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library axcelerator;
library techmap;
use techmap.axcomp.all;

entity grlfpw_0_axcelerator is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector (4 downto 0);
  cpi_d_pc : in std_logic_vector (31 downto 0);
  cpi_d_inst : in std_logic_vector (31 downto 0);
  cpi_d_cnt : in std_logic_vector (1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector (31 downto 0);
  cpi_a_inst : in std_logic_vector (31 downto 0);
  cpi_a_cnt : in std_logic_vector (1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector (31 downto 0);
  cpi_e_inst : in std_logic_vector (31 downto 0);
  cpi_e_cnt : in std_logic_vector (1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector (31 downto 0);
  cpi_m_inst : in std_logic_vector (31 downto 0);
  cpi_m_cnt : in std_logic_vector (1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector (31 downto 0);
  cpi_x_inst : in std_logic_vector (31 downto 0);
  cpi_x_cnt : in std_logic_vector (1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector (31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector (4 downto 0);
  cpi_dbg_data : in std_logic_vector (31 downto 0);
  cpo_data : out std_logic_vector (31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector (1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector (31 downto 0);
  rfi1_rd1addr : out std_logic_vector (3 downto 0);
  rfi1_rd2addr : out std_logic_vector (3 downto 0);
  rfi1_wraddr : out std_logic_vector (3 downto 0);
  rfi1_wrdata : out std_logic_vector (31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector (3 downto 0);
  rfi2_rd2addr : out std_logic_vector (3 downto 0);
  rfi2_wraddr : out std_logic_vector (3 downto 0);
  rfi2_wrdata : out std_logic_vector (31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector (31 downto 0);
  rfo1_data2 : in std_logic_vector (31 downto 0);
  rfo2_data1 : in std_logic_vector (31 downto 0);
  rfo2_data2 : in std_logic_vector (31 downto 0));
end grlfpw_0_axcelerator;

architecture beh of grlfpw_0_axcelerator is
  signal CPI_D_INST_0 : std_logic_vector (11 downto 9);
  signal CPI_DBG_ADDR_0 : std_logic_vector (0 to 0);
  signal CPI_DBG_ADDR_0_0 : std_logic_vector (0 to 0);
  signal CPI_DBG_ADDR_1 : std_logic_vector (0 to 0);
  signal CPI_DBG_ADDR_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_COMB_MEXC_1 : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_COMB_RS1_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_RS2_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_COMB_V_E_STDATA_1 : std_logic_vector (31 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_AEXC_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_CEXC_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_FCC_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_RD_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_TEM_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_I_INST_1 : std_logic_vector (31 downto 0);
  signal GRLFPC2_0_COMB_V_I_PC_1 : std_logic_vector (31 downto 2);
  signal GRLFPC2_0_COMB_V_I_RES_1 : std_logic_vector (63 downto 29);
  signal GRLFPC2_0_COMB_V_I_RES_6 : std_logic_vector (63 to 63);
  signal GRLFPC2_0_COMB_V_I_RES_6_CM8I : std_logic_vector (63 to 63);
  signal GRLFPC2_0_COMB_V_STATE_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_STATE_1_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_COMB_V_STATE_7 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_COMB_WRDATA_4 : std_logic_vector (62 downto 0);
  signal GRLFPC2_0_FPO_CC : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_FPO_EXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_FPO_EXP : std_logic_vector (10 downto 0);
  signal GRLFPC2_0_FPO_FRAC : std_logic_vector (54 downto 3);
  signal GRLFPC2_0_FPO_FRAC_0 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONCODES_1_CM8I : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4 : std_logic_vector (38 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I : std_logic_vector (50 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I : std_logic_vector (56 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N : std_logic_vector (57 downto 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N_CM8I : std_logic_vector (57 downto 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3 : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N : std_logic_vector (50 downto 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8 : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0 : std_logic_vector (57 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I : std_logic_vector (57 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_TZ : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_2 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_4 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I : std_logic_vector (55 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14 : std_logic_vector (142 to 142);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_CM8I : std_logic_vector (142 to 142);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23 : std_logic_vector (113 downto 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49 : std_logic_vector (258 to 258);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_50 : std_logic_vector (316 to 316);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1 : std_logic_vector (3 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2 : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_CM8I : std_logic_vector (3 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_N : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4 : std_logic_vector (57 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I : std_logic_vector (11 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8 : std_logic_vector (57 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I : std_logic_vector (57 downto 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_CM8I : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_2_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP : std_logic_vector (8 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0 : std_logic_vector (8 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0 : std_logic_vector (8 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1 : std_logic_vector (8 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0 : std_logic_vector (4 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2 : std_logic_vector (8 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3 : std_logic_vector (8 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4 : std_logic_vector (8 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5 : std_logic_vector (8 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6 : std_logic_vector (8 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7 : std_logic_vector (6 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8 : std_logic_vector (6 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9 : std_logic_vector (6 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10 : std_logic_vector (4 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_QUOBITS : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1 : std_logic_vector (55 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I : std_logic_vector (47 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N : std_logic_vector (57 downto 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8 : std_logic_vector (57 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I : std_logic_vector (57 downto 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N : std_logic_vector (54 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N_CM8I : std_logic_vector (49 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4_CM8I : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5_CM8I : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6_CM8I : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7_CM8I : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8_CM8I : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11_CM8I : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12_CM8I : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13_CM8I : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14_CM8I : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15_CM8I : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0_N : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17_0 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17_CM8I : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18_0 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19_0 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19_CM8I : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20_CM8I : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21_CM8I : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22_CM8I : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23_CM8I : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24_CM8I : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25_CM8I : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27_CM8I : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28_CM8I : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_0 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_CM8I : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31_CM8I : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32_CM8I : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33_CM8I : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34_CM8I : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35 : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35_CM8I : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36_CM8I : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37_0 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37_CM8I : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39_CM8I : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40_CM8I : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41_CM8I : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42_CM8I : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43_CM8I : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_0 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_CM8I : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45_CM8I : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47_CM8I : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48_0 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48_CM8I : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49_CM8I : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50_CM8I : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52_CM8I : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53_CM8I : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61_CM8I : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_CM8I : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63_CM8I : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64_CM8I : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66_0 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67_CM8I : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68_CM8I : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69_CM8I : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70_CM8I : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71_CM8I : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72_CM8I : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73_CM8I : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0_CM8I : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75_CM8I : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0_CM8I : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_77_0 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78_CM8I : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79_CM8I : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80_CM8I : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81_CM8I : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83_0 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84_CM8I : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85_CM8I : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87_CM8I : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88_0 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89_CM8I : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90_CM8I : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92_CM8I : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93_CM8I : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95_CM8I : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96_CM8I : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97_CM8I : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98_CM8I : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99_CM8I : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100_CM8I : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101_CM8I : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103_CM8I : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104_CM8I : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105_CM8I : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106_CM8I : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108_CM8I : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109_CM8I : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_110_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0_CM8I : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_CM8I : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119_CM8I : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_CM8I : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123_CM8I : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124_CM8I : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125_CM8I : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126_CM8I : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127_CM8I : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128_CM8I : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_CM8I : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_CM8I : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131_CM8I : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132_CM8I : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133_CM8I : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134_CM8I : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0_CM8I : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136_CM8I : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_CM8I : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139_CM8I : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_CM8I : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141_CM8I : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143_CM8I : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144_CM8I : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145_CM8I : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0_CM8I : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147 : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147_CM8I : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148_CM8I : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0_CM8I : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_0 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152_CM8I : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153_CM8I : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_CM8I : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155_CM8I : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156_CM8I : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157_CM8I : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159_CM8I : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160_CM8I : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161_CM8I : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162_CM8I : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164_CM8I : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165_CM8I : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_113_0 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_170 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_112_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_169 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_54 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_111 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_168 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53_CM8I : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_110 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_167 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52_CM8I : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_109 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_166 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_108 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_165 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50_CM8I : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_107 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ_CM8I : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_49 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_163 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_48 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ_CM8I : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_162 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_104 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_161 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_103 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_45 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_159 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44_CM8I : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_101 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158_CM8I : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_43 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ_CM8I : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_157 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_99 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_156 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_41 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_98 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_155 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_40 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_97 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_154 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_39 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_96 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_153 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_38 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_95 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_152 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_37 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_94 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_151 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_36 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_93 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_150 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35 : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35_CM8I : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_92 : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_149 : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34_CM8I : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_91 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_148 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_33 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N_CM8I : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_147 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_89 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_146 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_31 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_88 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_145 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_30 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_87 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_144 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_29 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_86 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_143 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_28 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ_CM8I : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_142 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ_CM8I : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_141 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_140 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_25_0 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_82 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_139 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_24 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81_CM8I : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_138 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_80 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_137 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_22 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_79 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_136 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_21 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_78 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_135 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_20 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_77 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_134 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_19 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_76 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_133 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_18 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_75 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_132 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17_CM8I : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_74 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_131 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_16 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_73 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_130 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15_CM8I : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_72 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_129 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14_CM8I : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_71 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_128 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_13 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_70 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_127 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_12 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_69 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_126 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_11 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_68 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_125 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_67 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_124 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_9 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_66 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_123 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_8 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_65 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_122 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_7 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_64 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_121 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_6 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_63 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_120 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_5 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_62 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_119 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_4 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_61 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118_CM8I : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_3 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ_CM8I : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_117 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_59 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_116 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS : std_logic_vector (12 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS : std_logic_vector (12 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I : std_logic_vector (12 downto 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS : std_logic_vector (56 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_CM8I : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I : std_logic_vector (56 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK : std_logic_vector (4 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_N : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_N_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_EXMIPTR : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_0_N_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I : std_logic_vector (7 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_2_0 : std_logic_vector (65 to 65);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14 : std_logic_vector (77 to 77);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0 : std_logic_vector (77 to 77);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_2 : std_logic_vector (77 to 77);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6 : std_logic_vector (3 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STATUS_1 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8 : std_logic_vector (9 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8_CM8I : std_logic_vector (9 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_10 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1 : std_logic_vector (9 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0_N : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4_N : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4_N_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_6 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_6_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_CM8I : std_logic_vector (5 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_A2_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_A7_0_N : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_O2_0_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0 : std_logic_vector (3 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_2 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A2_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_1_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_CM8I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1 : std_logic_vector (54 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19 : std_logic_vector (98 downto 84);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I : std_logic_vector (9 downto 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPRF_DOUT1_M : std_logic_vector (63 to 63);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE : std_logic_vector (12 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI : std_logic_vector (12 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19 : std_logic_vector (61 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0 : std_logic_vector (51 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0 : std_logic_vector (62 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I : std_logic_vector (59 downto 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1 : std_logic_vector (58 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_1 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I : std_logic_vector (58 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_TZ_TZ : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2 : std_logic_vector (55 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_CM8I : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_N : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_N_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_TZ : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3 : std_logic_vector (62 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I : std_logic_vector (62 downto 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_N : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_N_CM8I : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_TZ_N : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_TZ_N_CM8I : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4 : std_logic_vector (58 downto 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I : std_logic_vector (58 downto 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N : std_logic_vector (28 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N_CM8I : std_logic_vector (28 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5 : std_logic_vector (58 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I : std_logic_vector (31 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_N : std_logic_vector (62 to 62);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6 : std_logic_vector (62 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I : std_logic_vector (62 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_N : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_N_CM8I : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7 : std_logic_vector (59 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_CM8I : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N : std_logic_vector (32 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N_CM8I : std_logic_vector (32 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8 : std_logic_vector (59 downto 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I : std_logic_vector (59 downto 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N : std_logic_vector (58 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I : std_logic_vector (58 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_TZ : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_TZ_CM8I : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9 : std_logic_vector (59 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_0_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N : std_logic_vector (53 downto 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10 : std_logic_vector (57 downto 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I : std_logic_vector (52 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_N : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11 : std_logic_vector (57 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_CM8I : std_logic_vector (53 downto 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_N : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_N_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12 : std_logic_vector (55 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I : std_logic_vector (54 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N : std_logic_vector (59 downto 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N_CM8I : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13 : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14 : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_1 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I : std_logic_vector (57 downto 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_N : std_logic_vector (58 downto 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15 : std_logic_vector (58 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I : std_logic_vector (58 downto 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16 : std_logic_vector (58 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16_CM8I : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17 : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_CM8I : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_N : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_N_CM8I : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18 : std_logic_vector (55 downto 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_CM8I : std_logic_vector (55 downto 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_N : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_N_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19 : std_logic_vector (55 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_CM8I : std_logic_vector (55 downto 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_N : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_N_CM8I : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20 : std_logic_vector (57 downto 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21 : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I : std_logic_vector (59 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_CM8I : std_logic_vector (28 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_1_0 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_2_CM8I : std_logic_vector (28 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_CM8I : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_CM8I : std_logic_vector (28 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_0_0 : std_logic_vector (62 to 62);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_1_1 : std_logic_vector (62 to 62);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_5_1 : std_logic_vector (62 to 62);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_CM8I : std_logic_vector (62 to 62);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_1_N : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_0 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_1_N : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_12_0 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_0_0 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_CM8I : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_0 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_4_CM8I : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_13_1 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_0 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_0_CM8I : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_CM8I : std_logic_vector (53 downto 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_CM8I : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_0 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_6_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_CM8I : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_0 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_1 : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_11_1 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_17_1 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_CM8I : std_logic_vector (54 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_N_CM8I : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_1 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_0 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_CM8I : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_1_N : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_0 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_1 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_1 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_19_0 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_1_0_N : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_CM8I : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_N_CM8I : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_2_CM8I : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_3_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_1 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_5_CM8I : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_0 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_1 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_7_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_8_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_10_0 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_14_0 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_0 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_CM8I : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_0_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_1_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_3_CM8I : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_4_0 : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_5_0 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_0 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_1 : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_7_0 : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_1 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_10_1 : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_11_1 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_13_0 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_15_0 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_19_0 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_20_0_N : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_21_CM8I : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_22_1 : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_CM8I : std_logic_vector (59 to 59);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_0_0 : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_0 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_CM8I : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_0 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_1_N : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_1_N_CM8I : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_1 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_N_CM8I : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_1 : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_8_CM8I : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_11_0_N : std_logic_vector (58 to 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_15_0 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_17_1 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_19_0 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_CM8I : std_logic_vector (58 downto 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_1 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_N_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_1_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_2_1 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_3_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_4_1 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_5_CM8I : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_0_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_9_1 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_10_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_12_0 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_18_1 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_20_0 : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_21_0 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_23_1 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I : std_logic_vector (58 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I : std_logic_vector (57 downto 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N : std_logic_vector (43 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I : std_logic_vector (43 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_11_CM8I : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O28_CM8I : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1 : std_logic_vector (50 downto 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0 : std_logic_vector (7 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0_CM8I : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_1 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_2_N_CM8I : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I : std_logic_vector (50 downto 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N : std_logic_vector (30 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N_CM8I : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2 : std_logic_vector (61 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I : std_logic_vector (61 downto 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N : std_logic_vector (41 downto 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I : std_logic_vector (41 downto 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3 : std_logic_vector (61 downto 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I : std_logic_vector (38 downto 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_N : std_logic_vector (25 downto 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4 : std_logic_vector (51 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I : std_logic_vector (51 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_N : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_TZ : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5 : std_logic_vector (61 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_0 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_CM8I : std_logic_vector (7 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N : std_logic_vector (33 downto 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N_CM8I : std_logic_vector (33 downto 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6 : std_logic_vector (38 downto 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_CM8I : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N : std_logic_vector (26 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N_CM8I : std_logic_vector (26 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7 : std_logic_vector (51 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_0 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I : std_logic_vector (51 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N : std_logic_vector (61 downto 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N_CM8I : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8 : std_logic_vector (61 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I : std_logic_vector (61 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9 : std_logic_vector (61 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_CM8I : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N : std_logic_vector (50 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N_CM8I : std_logic_vector (50 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10 : std_logic_vector (51 downto 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_CM8I : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N : std_logic_vector (17 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N_CM8I : std_logic_vector (17 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11 : std_logic_vector (49 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_CM8I : std_logic_vector (36 downto 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_N : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12 : std_logic_vector (51 downto 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12_CM8I : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12_N : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13 : std_logic_vector (49 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13_CM8I : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N_CM8I : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N : std_logic_vector (51 downto 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N_CM8I : std_logic_vector (51 downto 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_16_N : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_16_N_CM8I : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_17 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_17_N : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_18 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_18_CM8I : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0 : std_logic_vector (42 downto 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_CM8I : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_N : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_0 : std_logic_vector (62 to 62);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0 : std_logic_vector (45 downto 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_0 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0 : std_logic_vector (36 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0 : std_logic_vector (50 downto 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_3_0 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_5_0 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0 : std_logic_vector (49 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_N_CM8I : std_logic_vector (49 downto 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I : std_logic_vector (61 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0 : std_logic_vector (56 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_TZ : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_TZ_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_1_N : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_1_N_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2 : std_logic_vector (60 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4 : std_logic_vector (60 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_5 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_5_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6 : std_logic_vector (60 downto 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_0 : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_CM8I : std_logic_vector (60 downto 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_8 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_8_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_9 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_9_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_10 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_10_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_11 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_11_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12 : std_logic_vector (60 downto 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_CM8I : std_logic_vector (60 downto 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_N : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_N_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13 : std_logic_vector (60 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14 : std_logic_vector (60 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I : std_logic_vector (56 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15 : std_logic_vector (56 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15_N : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15_N_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16 : std_logic_vector (56 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16_CM8I : std_logic_vector (47 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17 : std_logic_vector (56 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18 : std_logic_vector (56 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18_CM8I : std_logic_vector (56 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19 : std_logic_vector (56 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_N : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_N_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_20_N : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_20_N_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_21_N : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N : std_logic_vector (47 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N : std_logic_vector (56 downto 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_24_N : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_24_N_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_0_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_1_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_2_1 : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_2_CM8I : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_3_0 : std_logic_vector (60 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_7_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_8_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_9_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_10_0 : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_19_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_N_CM8I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_0_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_1_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_2_0 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_2_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_0 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_0_CM8I : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_4_0 : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_10_1 : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_23_0 : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_O28_2_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_M2_CM8I : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0 : std_logic_vector (38 downto 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0_0_CM8I : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_CM8I : std_logic_vector (26 downto 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_CM8I : std_logic_vector (36 downto 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I : std_logic_vector (50 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_1 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_21 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH : std_logic_vector (377 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0 : std_logic_vector (111 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0 : std_logic_vector (52 downto 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1 : std_logic_vector (54 to 54);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I : std_logic_vector (244 downto 232);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I : std_logic_vector (85 downto 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0 : std_logic_vector (83 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I : std_logic_vector (34 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11 : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12 : std_logic_vector (84 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13 : std_logic_vector (78 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL : std_logic_vector (16 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I : std_logic_vector (16 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_M : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_M_0_0 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH : std_logic_vector (375 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0 : std_logic_vector (375 downto 374);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I : std_logic_vector (375 downto 171);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1 : std_logic_vector (375 to 375);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I : std_logic_vector (112 downto 95);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I : std_logic_vector (115 downto 58);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_5_CM8I : std_logic_vector (55 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_7_CM8I : std_logic_vector (55 to 55);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I : std_logic_vector (244 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_D_CM8I : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_S_CM8I : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1 : std_logic_vector (54 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I : std_logic_vector (17 downto 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2 : std_logic_vector (56 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I : std_logic_vector (54 downto 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2 : std_logic_vector (50 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I : std_logic_vector (17 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N : std_logic_vector (49 downto 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N_CM8I : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SLCONTROL : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN : std_logic_vector (5 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_N : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_DIVMULTV : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_DIVMULTV_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI : std_logic_vector (7 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT : std_logic_vector (8 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_1_TZ : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN4_TEMP_U_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE : std_logic_vector (12 downto 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI : std_logic_vector (12 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI : std_logic_vector (57 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1 : std_logic_vector (68 to 68);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0 : std_logic_vector (68 to 68);
  signal GRLFPC2_0_OP1 : std_logic_vector (63 downto 32);
  signal GRLFPC2_0_OP2 : std_logic_vector (63 downto 32);
  signal GRLFPC2_0_R_A_RF1REN : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_R_A_RF2REN : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_R_A_RS1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_A_RS2 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_FSR_AEXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_FSR_CEXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_FSR_FTT : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_R_FSR_RD : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_R_FSR_TEM : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_I_CC : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_R_I_EXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_I_EXC_1_CM8I : std_logic_vector (2 to 2);
  signal GRLFPC2_0_R_I_INST : std_logic_vector (31 downto 0);
  signal GRLFPC2_0_R_I_PC : std_logic_vector (31 downto 2);
  signal GRLFPC2_0_R_I_RES : std_logic_vector (63 downto 0);
  signal GRLFPC2_0_R_STATE : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_RF1REN_CM8I : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_RF2REN_CM8I : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_V_FSR_FTT_1 : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_V_FSR_FTT_1_CM8I : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_WREN1_M : std_logic_vector (0 to 0);
  signal GRLFPC2_0_WREN1_M_CM8I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_WREN1_M_N : std_logic_vector (0 to 0);
  signal GRLFPC2_0_WREN210_M_N : std_logic_vector (340 to 340);
  signal NN_1 : std_logic ;
  signal NN_2 : std_logic ;
  signal N_1 : std_logic ;
  signal N_5577 : std_logic ;
  signal N_5579 : std_logic ;
  signal N_5580 : std_logic ;
  signal N_5581 : std_logic ;
  signal N_7971_N : std_logic ;
  signal N_7973 : std_logic ;
  signal N_7974 : std_logic ;
  signal N_7976 : std_logic ;
  signal N_7979 : std_logic ;
  signal N_7980 : std_logic ;
  signal N_7983 : std_logic ;
  signal N_7984 : std_logic ;
  signal N_7986 : std_logic ;
  signal N_7988 : std_logic ;
  signal N_7993 : std_logic ;
  signal N_8050 : std_logic ;
  signal NN_3 : std_logic ;
  signal NN_4 : std_logic ;
  signal CPI_DBG_ENABLE_0 : std_logic ;
  signal CPI_DBG_FSR_0 : std_logic ;
  signal CPI_DBG_FSR_0_0 : std_logic ;
  signal CPI_DBG_FSR_1 : std_logic ;
  signal CPI_DBG_FSR_2 : std_logic ;
  signal CPO_CC_0_INT_2 : std_logic ;
  signal CPO_CC_1_INT_3 : std_logic ;
  signal CPO_EXC_INT_1 : std_logic ;
  signal CPO_HOLDN_INT_4 : std_logic ;
  signal GRLFPC2_0_I_349_CM8I : std_logic ;
  signal GRLFPC2_0_I_352_1 : std_logic ;
  signal GRLFPC2_0_I_352_2 : std_logic ;
  signal GRLFPC2_0_I_352_4 : std_logic ;
  signal GRLFPC2_0_I_378_CM8I : std_logic ;
  signal GRLFPC2_0_I_388_CM8I : std_logic ;
  signal GRLFPC2_0_I_422_1_N_CM8I : std_logic ;
  signal GRLFPC2_0_I_422_CM8I : std_logic ;
  signal GRLFPC2_0_I_423_0 : std_logic ;
  signal GRLFPC2_0_I_423_0_CM8I : std_logic ;
  signal GRLFPC2_0_N_1 : std_logic ;
  signal GRLFPC2_0_N_12 : std_logic ;
  signal GRLFPC2_0_N_16_1 : std_logic ;
  signal GRLFPC2_0_N_17 : std_logic ;
  signal GRLFPC2_0_N_17_1 : std_logic ;
  signal GRLFPC2_0_N_161 : std_logic ;
  signal GRLFPC2_0_N_163 : std_logic ;
  signal GRLFPC2_0_N_164 : std_logic ;
  signal GRLFPC2_0_N_165 : std_logic ;
  signal GRLFPC2_0_N_166 : std_logic ;
  signal GRLFPC2_0_N_167 : std_logic ;
  signal GRLFPC2_0_N_169 : std_logic ;
  signal GRLFPC2_0_N_171 : std_logic ;
  signal GRLFPC2_0_N_173 : std_logic ;
  signal GRLFPC2_0_N_331 : std_logic ;
  signal GRLFPC2_0_N_335 : std_logic ;
  signal GRLFPC2_0_N_353_1 : std_logic ;
  signal GRLFPC2_0_N_548 : std_logic ;
  signal GRLFPC2_0_N_552 : std_logic ;
  signal GRLFPC2_0_N_640 : std_logic ;
  signal GRLFPC2_0_N_642 : std_logic ;
  signal GRLFPC2_0_N_643 : std_logic ;
  signal GRLFPC2_0_N_644 : std_logic ;
  signal GRLFPC2_0_N_645 : std_logic ;
  signal GRLFPC2_0_N_646 : std_logic ;
  signal GRLFPC2_0_N_647 : std_logic ;
  signal GRLFPC2_0_N_655 : std_logic ;
  signal GRLFPC2_0_N_656 : std_logic ;
  signal GRLFPC2_0_N_658 : std_logic ;
  signal GRLFPC2_0_N_659 : std_logic ;
  signal GRLFPC2_0_N_664 : std_logic ;
  signal GRLFPC2_0_N_665 : std_logic ;
  signal GRLFPC2_0_N_666 : std_logic ;
  signal GRLFPC2_0_N_667 : std_logic ;
  signal GRLFPC2_0_N_668 : std_logic ;
  signal GRLFPC2_0_N_816 : std_logic ;
  signal GRLFPC2_0_N_817 : std_logic ;
  signal GRLFPC2_0_N_818 : std_logic ;
  signal GRLFPC2_0_N_819 : std_logic ;
  signal GRLFPC2_0_N_820 : std_logic ;
  signal GRLFPC2_0_N_849 : std_logic ;
  signal GRLFPC2_0_N_857 : std_logic ;
  signal GRLFPC2_0_N_865 : std_logic ;
  signal GRLFPC2_0_N_866 : std_logic ;
  signal GRLFPC2_0_N_878 : std_logic ;
  signal GRLFPC2_0_N_879 : std_logic ;
  signal GRLFPC2_0_N_880 : std_logic ;
  signal GRLFPC2_0_N_881 : std_logic ;
  signal GRLFPC2_0_N_882 : std_logic ;
  signal GRLFPC2_0_N_895 : std_logic ;
  signal GRLFPC2_0_N_897 : std_logic ;
  signal GRLFPC2_0_N_898 : std_logic ;
  signal GRLFPC2_0_N_900 : std_logic ;
  signal GRLFPC2_0_N_901 : std_logic ;
  signal GRLFPC2_0_N_902 : std_logic ;
  signal GRLFPC2_0_N_903 : std_logic ;
  signal GRLFPC2_0_N_904 : std_logic ;
  signal GRLFPC2_0_N_905 : std_logic ;
  signal GRLFPC2_0_N_906 : std_logic ;
  signal GRLFPC2_0_N_907 : std_logic ;
  signal GRLFPC2_0_N_908 : std_logic ;
  signal GRLFPC2_0_N_909 : std_logic ;
  signal GRLFPC2_0_N_910 : std_logic ;
  signal GRLFPC2_0_N_911 : std_logic ;
  signal GRLFPC2_0_N_912 : std_logic ;
  signal GRLFPC2_0_N_913 : std_logic ;
  signal GRLFPC2_0_N_914 : std_logic ;
  signal GRLFPC2_0_N_915 : std_logic ;
  signal GRLFPC2_0_N_916 : std_logic ;
  signal GRLFPC2_0_N_917 : std_logic ;
  signal GRLFPC2_0_N_918 : std_logic ;
  signal GRLFPC2_0_N_919 : std_logic ;
  signal GRLFPC2_0_N_920 : std_logic ;
  signal GRLFPC2_0_N_923 : std_logic ;
  signal GRLFPC2_0_N_924 : std_logic ;
  signal GRLFPC2_0_N_925 : std_logic ;
  signal GRLFPC2_0_N_926 : std_logic ;
  signal GRLFPC2_0_N_927 : std_logic ;
  signal GRLFPC2_0_N_929 : std_logic ;
  signal GRLFPC2_0_N_932 : std_logic ;
  signal GRLFPC2_0_N_954 : std_logic ;
  signal GRLFPC2_0_N_1058 : std_logic ;
  signal GRLFPC2_0_N_1059 : std_logic ;
  signal GRLFPC2_0_N_1063 : std_logic ;
  signal GRLFPC2_0_N_1063_3 : std_logic ;
  signal GRLFPC2_0_N_1080 : std_logic ;
  signal GRLFPC2_0_N_1093 : std_logic ;
  signal GRLFPC2_0_N_1104 : std_logic ;
  signal GRLFPC2_0_N_1105 : std_logic ;
  signal GRLFPC2_0_N_1108 : std_logic ;
  signal GRLFPC2_0_N_1109_N : std_logic ;
  signal GRLFPC2_0_N_1123 : std_logic ;
  signal GRLFPC2_0_N_1127 : std_logic ;
  signal GRLFPC2_0_N_1132 : std_logic ;
  signal GRLFPC2_0_N_1132_1_N : std_logic ;
  signal GRLFPC2_0_N_1133 : std_logic ;
  signal GRLFPC2_0_ANNULRES_0_SQMUXA_3_1 : std_logic ;
  signal GRLFPC2_0_ANNULRES_0_SQMUXA_4_1 : std_logic ;
  signal GRLFPC2_0_ANNULRES_1_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0 : std_logic ;
  signal GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_ANNULFPU_1 : std_logic ;
  signal GRLFPC2_0_COMB_ANNULFPU_1_U_0 : std_logic ;
  signal GRLFPC2_0_COMB_ANNULRES_1 : std_logic ;
  signal GRLFPC2_0_COMB_CCWR4_1 : std_logic ;
  signal GRLFPC2_0_COMB_CCWR4_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_CCWR4_1_0_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ3 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ3_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ6_N : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ6_N_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ12 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ13 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV2 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV2_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV2_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV4_2 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV4_3 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV5 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV5_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV6 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV7 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV7_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV11 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV12 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_RS2D5 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_RS2D5_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_RS2D5_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_ST : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_ST_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_3 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_4 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_5 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_WREN210 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN3_OP : std_logic ;
  signal GRLFPC2_0_COMB_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_ISFPOP2_1 : std_logic ;
  signal GRLFPC2_0_COMB_ISFPOP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_LOCK_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_DEPCHECK : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_DEPCHECK_1 : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_1 : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_UN6_DEPCHECK : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_UN8_DEPCHECK : std_logic ;
  signal GRLFPC2_0_COMB_QNE2 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_1 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_1_1 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_0 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_0_0 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_1 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_2 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_3 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_4 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_5 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3_6 : std_logic ;
  signal GRLFPC2_0_COMB_RS1D_1 : std_logic ;
  signal GRLFPC2_0_COMB_RS1V_1_I_A4_0_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_RS1V_1_I_A4_0_1_1 : std_logic ;
  signal GRLFPC2_0_COMB_RS2_1_SN_N_2 : std_logic ;
  signal GRLFPC2_0_COMB_RS2_1_SN_N_2_0 : std_logic ;
  signal GRLFPC2_0_COMB_RS2D_1 : std_logic ;
  signal GRLFPC2_0_COMB_RSDECODE_UN1_FPCI : std_logic ;
  signal GRLFPC2_0_COMB_SEQERR_UN7_OP : std_logic ;
  signal GRLFPC2_0_COMB_SEQERR_UN7_OP_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_SEQERR_UN11_OP_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_2 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_3 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_0_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_2 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_2_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_4_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN1_MEXC : std_logic ;
  signal GRLFPC2_0_COMB_UN1_MEXC_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_MEXC_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN1_R_A_RS1_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_R_A_RS1_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_R_A_RS1_1_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_R_A_RS1_1_2 : std_logic ;
  signal GRLFPC2_0_COMB_UN2_HOLDN : std_logic ;
  signal GRLFPC2_0_COMB_UN2_HOLDN_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN2_HOLDN_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN2_HOLDN_2 : std_logic ;
  signal GRLFPC2_0_COMB_UN2_HOLDN_3 : std_logic ;
  signal GRLFPC2_0_COMB_UN3_HOLDN : std_logic ;
  signal GRLFPC2_0_COMB_UN3_HOLDN_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN4_LOCK : std_logic ;
  signal GRLFPC2_0_COMB_UN4_LOCK_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC_0_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC_2 : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC_3 : std_logic ;
  signal GRLFPC2_0_COMB_UN8_CCV_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN8_CCV_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_UN9_CCV : std_logic ;
  signal GRLFPC2_0_COMB_UN10_IUEXEC : std_logic ;
  signal GRLFPC2_0_COMB_UN10_IUEXEC_0 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFQ_1_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFQ_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_LD_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_LD_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_V_A_SEQERR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_ST_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_LD_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_STDATA2 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_STDATA2_0 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_STDATA2_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_STDATA2_2 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_NONSTD_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3 : std_logic ;
  signal GRLFPC2_0_COMB_V_I_EXEC_4 : std_logic ;
  signal GRLFPC2_0_COMB_V_I_EXEC_4_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_V_I_V6 : std_logic ;
  signal GRLFPC2_0_COMB_V_I_V_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_I_V_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_V_M_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_M_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_M_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_M_LD_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_MK_LDOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_MK_RST_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_MK_RST_1_3 : std_logic ;
  signal GRLFPC2_0_COMB_V_STATE12 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_LD_1 : std_logic ;
  signal GRLFPC2_0_COMB_WREN1_1_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_WREN1_9 : std_logic ;
  signal GRLFPC2_0_COMB_WREN1_9_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_WREN2_9 : std_logic ;
  signal GRLFPC2_0_COMB_WREN2_9S_IV_CM8I : std_logic ;
  signal GRLFPC2_0_COMB_WREN22 : std_logic ;
  signal GRLFPC2_0_COMB_WRRES4 : std_logic ;
  signal GRLFPC2_0_COMB_WRRES4_0 : std_logic ;
  signal GRLFPC2_0_FPI_LDOP : std_logic ;
  signal GRLFPC2_0_FPI_LDOP_0 : std_logic ;
  signal GRLFPC2_0_FPI_LDOP_1 : std_logic ;
  signal GRLFPC2_0_FPI_LDOP_2 : std_logic ;
  signal GRLFPC2_0_FPI_LDOP_3 : std_logic ;
  signal GRLFPC2_0_FPI_START : std_logic ;
  signal GRLFPC2_0_FPO_SIGN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1766_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1768_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1769_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1770_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1773_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1786_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1787_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1789_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1791_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1792_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1795_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1797_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1799_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1800_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1802_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1804_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1806_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1807_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1808_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1811_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1815_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1816_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1821_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1823_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1824_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1828_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1830_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1836_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1838_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_38 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_39 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_40 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_41 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_42 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_43 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_44 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_45 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_46 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_47 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_48 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_49 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_50 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_51 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_52 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_54 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_55 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_58 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_59 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_60 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_61 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_62 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_63 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_64 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_65 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_66 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_68 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_72 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_73 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_74 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_76 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_77 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_78 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_79 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_82 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_83 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_84 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_85 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_87 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_88 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_89 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_90 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_91 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_93 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_94 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_95 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_96 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_97 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_98 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_99 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_100 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_101 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_102 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_103 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_104 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_105 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_106 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_107 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_108 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_110 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_111 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_112 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_114 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_115 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_118 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_120 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_121 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_122 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_123 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_125 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_126 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_127 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_128 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_129 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_130 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_132 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_134 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_135 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_136 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_138 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_139 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_140 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_141 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_243 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_245_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_248 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_253 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_254 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_256 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_265 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_266 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_269 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_270 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_275 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_276 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_440_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_464 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_478_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_482 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_500 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_501 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_507 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_559 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_589 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_590 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_611 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_614 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_621 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_627 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_646 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_663 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_667_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_674_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_675 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_678 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_690 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_691_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_761 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_765 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_768 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_773 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_914 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_922 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_989 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_992 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_993 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_997 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1003 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1010 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1014 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1018_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1025 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1027 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1029 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1045_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1077 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1084 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1092 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1093 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1097 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1100 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1101 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1103_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1104 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1107 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1108 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1109_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1110_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1111 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1113 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1116 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1117 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1128 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1132 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1133 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1135 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1141 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1148 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1151 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1194 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1195 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1197 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1211 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1243 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1244 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1245 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1247 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1256 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1257 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1262 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1276 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1298_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1300 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1302 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1304 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1306 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1310 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1311_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1312 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1315 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1317 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1324 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1344 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1346 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1349 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1352 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1371 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1372 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1389_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1391 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1414 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1418 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1444 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1445 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1448 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1450 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1471 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1477 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1480 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1485 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1486 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1493 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1500 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1502_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1517 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1523 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1539 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1543 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1566 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1572 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1582 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1588 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1591_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1592 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1600 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1601 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1605 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1607 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1609 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1637 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1639 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1641 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1643 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1647 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1650 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1656 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1664 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1666 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2024_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2025 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2034 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2035 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2036 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2037 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2038 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2039 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2040 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2041 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2046 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2047 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2048 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2049 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2051 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2063 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2064 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2065 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2066 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2067 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2068 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2069 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2070 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2071 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2072 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2073 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2074 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2075 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2076 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2077 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2078 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2079 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2080 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2081 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2082 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2083 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2084 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2085 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2086 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2087 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2088 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2089 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2090 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2091 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2092 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2093 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2094 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2117 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2118 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2120 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2123 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2125 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2126 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2154 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2155 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2156 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2157 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2158 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2159 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2160 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2161 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2162 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2163 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2164 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2165 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2166 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2167 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2168 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2169 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2170 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2171 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2172 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2173 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2174 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2175 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2176 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2178 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2187 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2188 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2189 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2190 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2191 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2192 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2193 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2194 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2198 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2201 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2202 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2203 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2204 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2205 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2206 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2208 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2209 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2210 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2211 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2212 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2213 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2214 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2215 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2216 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2217 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2218 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2219 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2220 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2221 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2222 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2223 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2224 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2225 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2226 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2228 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2229 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2230 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2231 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2232 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2233 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2234 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2347 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2353 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2361 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2362 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2363 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2364 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2365 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2366 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2367 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2368 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2369 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2370 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2372 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2373 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2374 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2375 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2376 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2377 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2378 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2379 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2380 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2381 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2382 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2383 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2384 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2385 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2386 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2387 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2388 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2389 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2390 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2391 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2392 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2393 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2394 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2395 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2396 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2397 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2398 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2399 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2400 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2401 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2402 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2403 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2404 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2405 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2406 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2407 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2408 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2409 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2410 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2411 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2412 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2413 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2414 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2416 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2419 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2420_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2421_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2422_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2423_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2424_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2425_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2426_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2427_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2428_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2429_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2430_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2431_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2432_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2433_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2434_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2435_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2436_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2437_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2438_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2439_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2440_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2441_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2442_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2443_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2444_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2445_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2446_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2447_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2448_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2449_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2450_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2451_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2452_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2453_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2454_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2455_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2456_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2457_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2458_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2459_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2460_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2461_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2462_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2463_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2464_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2465_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2466_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2467 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2468_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2469_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2470_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2471_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2472_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2473 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2474_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2475 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2476 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2478 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2479 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2480 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2481 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2482 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2483 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2484 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2485 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2486 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2487 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2488 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2489 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2490 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2491 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2492 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2493 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2494 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2495 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2496 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2497 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2498 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2499 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2500 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2501 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2502 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2503 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2504 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2505 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2506 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2507 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2508 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2509 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2510 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2511 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2512 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2513 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2514 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2515 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2516 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2517 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2518 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2519 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2520 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2521 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2522 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2523 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2524 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2525 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2526 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2527 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2528 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2529 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2530 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2531 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2532 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2533 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2534 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2535 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2662 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2664 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2665 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2668 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2671 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2673 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2675 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2678 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2679 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2681 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2689 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2690 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2691 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2692 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2693 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2694 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2695 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2696 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2697 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2698 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2699 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2700 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2701 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2702 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2703 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2704 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2705 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2706 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2707 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2708 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2709 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2710 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2711 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2712 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2713 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2714 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2715 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2716 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2717 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2718 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2719 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2720 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2744 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2745 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2746 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2751 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2752 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2753 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2754 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2755 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2756 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2757 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2758 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2759 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2760 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2761 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2762 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2763 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2764 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2766 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2767 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2768 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2780 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2781 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2782 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2783 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2784 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2785 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2786 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2787 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2788 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2789 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2790 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2791 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2792 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2793 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2794 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2795 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2796 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2797 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2798 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2799 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2800 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2801 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2802 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2868 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2869 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2870 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2871 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2872 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2873 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2874 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2875 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2876 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2877 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2878 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2879 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2880 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2881 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2882 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2883 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2884 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2885 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2886 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2887 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2888 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2889 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2890 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2891 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2892 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2893 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2894 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2895 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2896 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2897 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2898 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2899 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2900 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2901 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2902 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2903 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2904 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2905 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2906 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2907 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2908 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2909 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2910 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2911 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2912 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2913 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2914 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2915 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2916 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2917 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2918 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2919 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2920 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2921 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2922 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2923 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2924 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2925 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2994 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2995 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2996 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2997 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2998 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2999 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3000 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3001 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3002 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3003 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3004 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3005 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3006 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3008 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3009 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3010 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3011 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3012 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3013 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3014 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3015 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3016 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3019 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3020 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3023 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3024 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3025 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3026 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3027 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3028 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3029 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3030 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3031 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3045 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3046 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3067 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3079 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3080 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3109 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3110 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3199 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3200 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3201 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3202 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3203 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3204 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3205 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3206 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3209 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3210 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3211 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3212 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3213 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3214 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3215 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3216 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3217 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3218 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3219 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3220 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3221 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3275_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3277 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3278 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3279 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3282 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3286 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3288 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3295 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3298 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3310_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3312 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3313_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3314_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3316_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3318 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3319 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3322_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3324 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3325 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3326 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3327 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3329 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3330 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3331 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3333 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3334_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3335_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3338_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3340 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3342 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3343 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3346 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3347 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3348 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3350 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3351 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3355_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3356 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3357_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3360 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3363_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3365_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3378 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3379 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3380 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3381 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3382 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3383 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3384 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3385 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3386 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3387 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3388 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3389 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3390 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3391 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3392 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3393 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3394 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3395 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3396 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3397 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3398 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3399 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3400 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3401 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3402 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3403 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3404 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3405 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3406 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3407 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3408 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3409 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3410 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3411 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3412 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3413 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3414 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3415 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3416 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3417 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3418 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3419 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3420 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3421 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3422 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3423 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3424 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3425 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3426 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3427 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3428 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3429 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3430 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3431 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3432 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3434_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3439_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3442_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3443_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3447_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3452_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3459_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3462_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3467_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3468_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3469_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3475_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3478_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3481_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3482_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3484_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3489_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3548 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3550_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3552 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3554 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3555 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3556 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3557 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3558_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3559_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3560_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3561 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3562_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3563 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3564_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3565 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3566_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3567_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3572 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3573 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3575_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3576_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3577_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3579_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3580 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3581_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3583_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3586_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3587_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3588_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3589_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3590 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3591_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3592 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3593 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3594_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3595_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3596_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3597 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3598_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3599_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3600_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3601_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3602_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3603_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3668 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3671 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3678 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3681 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3713 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3714 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3715 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3716 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3717 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3718 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3923_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3926 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3931 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3935 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3936 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3937 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3938 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3945 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3965_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3968 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3969 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3979 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3981 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3983 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3984 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3985_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3987 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3988 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3989 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3990 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3991 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3992 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4018 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4026 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4032 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4040 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4041 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4043 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4045 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4046 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4052 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4053 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4055_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4056 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4058 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4061 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4081 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4099 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4111_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4113 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4115_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4116 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4117 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4118 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4122 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4123 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4124_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4125_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4126 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4127_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4129_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4133 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4134 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4171 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4176_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4179 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4181 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4182_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4184_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4210 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4224 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4225 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4226 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4227_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4228 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4231_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4235 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4237 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4237_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4239 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4242 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4245 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4246 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4247 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4260 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4269 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4285 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4289 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4292 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4302 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4303 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4304 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4306 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4311 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4314 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4316 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4319 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4321 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4324 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4347 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4370 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4371 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4373 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4374 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4375_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4377 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4382 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4395 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4396 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4398 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4402 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4408_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4409 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4410 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4412 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4417 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4421 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4428_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4430 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4443 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4449 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4455_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4458 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4460 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4462 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4465 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4467 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4470_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4471 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4480 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4502 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4513_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4520 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4522 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4525_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4528_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4530 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4531 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4533 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4535 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4536 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4537 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4538 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4540 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4541 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4543 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4545_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4564 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4569_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4592 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4594 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4595 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4596 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4598_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4599_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4601 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4602 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4603 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4605 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4606 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4609 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4610 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4610_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4612 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4615 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4616_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4618_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4620 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4649_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4674 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4675 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4677 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4678_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4679 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4680 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4681 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4683 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4685 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4686 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4687_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4691 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4699 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4708 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4710 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4719 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4739 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4744 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4747 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4748_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4749 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4750 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4751 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4752 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4753 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4755 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4756_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4757 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4758 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4759 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4760 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4761 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4763 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4765 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4766_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4769 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4784 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4802 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4810 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4811 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4817 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4819 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4820 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4822 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4823_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4824 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4825 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4828 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4829 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4830 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4831 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4832 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4835 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4885_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4886 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4887_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4889_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4890_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4892_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4893 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4896 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4899 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4904 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4938 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4939_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4955 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4959 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4960 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4961 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4962_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4963 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4964 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4966_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4967 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4969 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4972 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4975 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4977_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4978_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4979 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4981 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5004 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5016_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5024 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5028 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5030 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5036 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5038 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5039 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5040 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5042 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5044 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5045 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5046 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5048 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5051_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5054 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5055_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5057 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5062 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5091 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5097_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5101_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5107 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5110 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5122 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5124 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5127 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5131 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5132_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5133 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5134 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5136 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5137 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5139 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5141_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5164 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5165 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5169 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5179 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5182 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5193_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5201 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5204 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5205 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5206 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5207 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5208_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5212 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5214 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5215 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5218 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5222_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5223_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5246 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5270 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5271 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5272 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5273 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5276 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5279_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5282 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5284_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5285 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5287 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5289 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5290 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5292 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5302 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5321_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5326 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5336_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5337 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5338 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5339_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5342 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5343 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5344 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5346 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5348_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5350_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5353 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5357 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5390 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5393 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5402 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5403 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5405_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5406 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5407 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5410 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5413 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5418 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_6545 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_6546 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SIGNRESULT_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTBINFNAN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_6_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_4_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN8_INFORCREGSN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN10_STKGEN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_STKOUT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN25_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN47_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN56_GEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTDIVISORBIT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN10_SHDVAR : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN28_SHDVAR : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN54_SHDVAR_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN54_SHDVAR_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN5_DIVMULTV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN86_DIVMULTV_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN111_DIVMULTV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN339_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN392_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN681_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN165_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN336_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN507_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN678_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN784_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN162_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN333_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN504_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN675_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN330_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN672_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN156_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN498_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN669_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN324_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN495_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN666_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN150_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN321_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN492_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN663_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN489_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN660_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN144_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN315_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN486_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN657_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN483_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN654_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN138_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN309_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN480_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN651_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN477_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN648_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN132_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN303_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN474_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN645_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN300_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN471_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN642_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN126_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN297_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN468_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN639_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN123_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN294_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN465_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN636_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN120_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN291_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN462_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN633_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN288_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN459_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN630_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN114_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN285_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN456_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN627_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN111_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN282_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN453_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN624_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN108_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN279_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN450_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN621_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN105_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN447_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN618_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN273_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN444_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN615_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN99_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN270_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN441_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN612_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN267_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN609_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN93_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN264_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN435_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN606_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN90_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN261_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN432_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN603_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN87_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN258_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN429_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN600_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN84_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN255_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN426_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN597_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN81_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN252_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN423_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN594_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN78_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN249_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN420_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN591_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN246_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN417_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN574_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN588_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN72_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN170_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN243_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN585_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN411_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN582_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN66_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN237_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN408_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN579_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN63_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN234_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN405_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN576_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN231_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN402_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN573_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN57_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN228_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN399_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN570_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN225_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN396_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN567_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN51_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN222_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN564_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN48_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN219_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN390_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN561_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN216_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN387_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN558_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN42_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN213_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN384_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN555_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN39_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN210_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN381_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN552_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN207_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN378_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN549_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN33_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN204_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN375_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN546_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN30_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN201_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN372_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN543_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN27_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN198_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN369_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN540_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN24_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN366_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN537_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN21_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN192_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN363_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN534_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN189_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN360_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN531_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN15_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN186_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN357_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN528_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN12_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN183_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN354_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN525_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN180_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN351_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN522_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN6_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN177_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN348_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN519_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN345_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN516_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN171_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN342_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN513_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_0_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN5_S_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_14_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_6_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_6_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_STICKYFORSR1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_NOTXZYFROMD : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN26_NOTXZYFROMD : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_34 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42_S : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42_S_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_48 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_55 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_2_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_3_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_4_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_5_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_0_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_15_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_16 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_16_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_21 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_22_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_25_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_26 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_27 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_27_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_4_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_6_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_7_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_10_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_13_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_21_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_23_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_0_D_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_0_S_2_N_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_SN_N_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN4_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN4_LOCUV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_3_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN21_LOCOV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN31_LOCOV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN4_NOTRESETORUNIMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN7_U_RDN_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN1_GRFPUS : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN5_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN10_AREGSIGN_SEL_M : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN2_SIGTAF38_37 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN58_SCTRL_NEW : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN5_NOTSHIFTCOUNT1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS_N : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_UN2_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_0_SQMUXA_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_N_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_7_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M5_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_S : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M6_0_CM8I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_AREGSIGN_SEL_INV_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_N_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_1 : std_logic ;
  signal NN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_N_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_N_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3 : std_logic ;
  signal GRLFPC2_0_M7_0 : std_logic ;
  signal GRLFPC2_0_M7_0_CM8I : std_logic ;
  signal GRLFPC2_0_MOV_5_SQMUXA : std_logic ;
  signal GRLFPC2_0_MOV_7_SQMUXA : std_logic ;
  signal GRLFPC2_0_R_A_AFQ : std_logic ;
  signal GRLFPC2_0_R_A_AFQ_0 : std_logic ;
  signal GRLFPC2_0_R_A_AFQ_1 : std_logic ;
  signal GRLFPC2_0_R_A_AFQ_2 : std_logic ;
  signal GRLFPC2_0_R_A_AFSR : std_logic ;
  signal GRLFPC2_0_R_A_AFSR_0 : std_logic ;
  signal GRLFPC2_0_R_A_AFSR_1 : std_logic ;
  signal GRLFPC2_0_R_A_AFSR_2 : std_logic ;
  signal GRLFPC2_0_R_A_FPOP : std_logic ;
  signal GRLFPC2_0_R_A_FPOP_0 : std_logic ;
  signal GRLFPC2_0_R_A_LD : std_logic ;
  signal GRLFPC2_0_R_A_MOV : std_logic ;
  signal GRLFPC2_0_R_A_RDD : std_logic ;
  signal GRLFPC2_0_R_A_RS1D : std_logic ;
  signal GRLFPC2_0_R_A_RS2D : std_logic ;
  signal GRLFPC2_0_R_A_SEQERR : std_logic ;
  signal GRLFPC2_0_R_A_ST : std_logic ;
  signal GRLFPC2_0_R_E_AFQ : std_logic ;
  signal GRLFPC2_0_R_E_AFSR : std_logic ;
  signal GRLFPC2_0_R_E_FPOP : std_logic ;
  signal GRLFPC2_0_R_E_LD : std_logic ;
  signal GRLFPC2_0_R_E_RDD : std_logic ;
  signal GRLFPC2_0_R_E_SEQERR : std_logic ;
  signal GRLFPC2_0_R_FSR_NONSTD : std_logic ;
  signal GRLFPC2_0_R_I_EXEC : std_logic ;
  signal GRLFPC2_0_R_I_RDD : std_logic ;
  signal GRLFPC2_0_R_I_V : std_logic ;
  signal GRLFPC2_0_R_M_AFQ : std_logic ;
  signal GRLFPC2_0_R_M_AFSR : std_logic ;
  signal GRLFPC2_0_R_M_FPOP : std_logic ;
  signal GRLFPC2_0_R_M_LD : std_logic ;
  signal GRLFPC2_0_R_M_RDD : std_logic ;
  signal GRLFPC2_0_R_M_SEQERR : std_logic ;
  signal GRLFPC2_0_R_MK_BUSY : std_logic ;
  signal GRLFPC2_0_R_MK_BUSY2 : std_logic ;
  signal GRLFPC2_0_R_MK_BUSY_0_2 : std_logic ;
  signal GRLFPC2_0_R_MK_HOLDN1 : std_logic ;
  signal GRLFPC2_0_R_MK_HOLDN2 : std_logic ;
  signal GRLFPC2_0_R_MK_LDOP : std_logic ;
  signal GRLFPC2_0_R_MK_RST : std_logic ;
  signal GRLFPC2_0_R_MK_RST2 : std_logic ;
  signal GRLFPC2_0_R_X_AFQ : std_logic ;
  signal GRLFPC2_0_R_X_AFSR : std_logic ;
  signal GRLFPC2_0_R_X_FPOP : std_logic ;
  signal GRLFPC2_0_R_X_FPOP_0 : std_logic ;
  signal GRLFPC2_0_R_X_LD : std_logic ;
  signal GRLFPC2_0_R_X_LD_0 : std_logic ;
  signal GRLFPC2_0_R_X_RDD : std_logic ;
  signal GRLFPC2_0_R_X_SEQERR : std_logic ;
  signal GRLFPC2_0_RS1D_CNST : std_logic ;
  signal GRLFPC2_0_RS1D_CNST_0_A2_0 : std_logic ;
  signal GRLFPC2_0_RS1D_CNST_0_A3_0_0_N : std_logic ;
  signal GRLFPC2_0_RS1D_CNST_0_O2_CM8I : std_logic ;
  signal GRLFPC2_0_RS1V10 : std_logic ;
  signal GRLFPC2_0_RS1V_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_RS2_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_UN1_FPCI_2_N : std_logic ;
  signal GRLFPC2_0_UN1_FPCI_2_N_CM8I : std_logic ;
  signal GRLFPC2_0_UN1_FPCI_3_0 : std_logic ;
  signal GRLFPC2_0_UN1_FPCI_3_1 : std_logic ;
  signal GRLFPC2_0_UN1_HOLDN_1 : std_logic ;
  signal GRLFPC2_0_UN1_HOLDN_1_0 : std_logic ;
  signal GRLFPC2_0_UN1_HOLDN_1_1 : std_logic ;
  signal GRLFPC2_0_UN1_HOLDN_1_2 : std_logic ;
  signal GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0 : std_logic ;
  signal GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0_CM8I : std_logic ;
  signal GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_1 : std_logic ;
  signal GRLFPC2_0_UN1_WREN1_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_UN1_WREN1_0_SQMUXA_CM8I : std_logic ;
  signal GRLFPC2_0_V_FSR_FTT_0_SQMUXA_2_1 : std_logic ;
  signal GRLFPC2_0_V_FSR_FTT_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0 : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0 : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_0 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_3 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_4 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_5 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA_6 : std_logic ;
  signal GRLFPC2_0_V_I_V_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_STATE_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_STATE_1_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_V_STATE_1_SQMUXA_CM8I : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_0 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_0_0 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_0 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_1 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_2 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_3 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_4 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_5 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1_6 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_3 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_4 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_5 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_6 : std_logic ;
  signal GRLFPC2_0_WRADDR_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_WREN1_0_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_WREN1_0_SQMUXA_3 : std_logic ;
  signal GRLFPC2_0_WREN2_2_SQMUXA_0 : std_logic ;
  signal HOLDN_0 : std_logic ;
  signal HOLDN_1 : std_logic ;
  signal HOLDN_I : std_logic ;
  signal HOLDN_I_0 : std_logic ;
  signal HOLDN_I_0_0 : std_logic ;
  signal HOLDN_I_0_1 : std_logic ;
  signal HOLDN_I_1 : std_logic ;
  signal HOLDN_I_1_0 : std_logic ;
  signal HOLDN_I_2 : std_logic ;
  signal HOLDN_I_3 : std_logic ;
  signal HOLDN_I_4 : std_logic ;
  signal HOLDN_I_5 : std_logic ;
  signal HOLDN_I_6 : std_logic ;
  signal HOLDN_I_7 : std_logic ;
  signal HOLDN_I_8 : std_logic ;
  signal HOLDN_I_9 : std_logic ;
  signal HOLDN_I_10 : std_logic ;
  signal HOLDN_I_11 : std_logic ;
  signal HOLDN_I_12 : std_logic ;
  signal HOLDN_I_13 : std_logic ;
  signal HOLDN_I_14 : std_logic ;
  signal HOLDN_I_15 : std_logic ;
  signal HOLDN_I_16 : std_logic ;
  signal HOLDN_I_17 : std_logic ;
  signal RFI1_WRDATA_31_INT_17 : std_logic ;
  signal RFI2_RD1ADDR_0_INT_5_INT_18 : std_logic ;
  signal RFI2_RD1ADDR_1_INT_6_INT_19 : std_logic ;
  signal RFI2_RD1ADDR_2_INT_7_INT_20 : std_logic ;
  signal RFI2_RD1ADDR_3_INT_8_INT_21 : std_logic ;
  signal RFI2_RD2ADDR_0_INT_9_INT_22 : std_logic ;
  signal RFI2_RD2ADDR_1_INT_10_INT_23 : std_logic ;
  signal RFI2_RD2ADDR_2_INT_11_INT_24 : std_logic ;
  signal RFI2_RD2ADDR_3_INT_12_INT_25 : std_logic ;
  signal RFI2_WRADDR_0_INT_13_INT_26 : std_logic ;
  signal RFI2_WRADDR_1_INT_14_INT_27 : std_logic ;
  signal RFI2_WRADDR_2_INT_15_INT_28 : std_logic ;
  signal RFI2_WRADDR_3_INT_16_INT_29 : std_logic ;
  signal RST_I : std_logic ;
begin
  NN_1 <= '0';
  x_GND_Z9619: GND port map (
      Y => NN_2);
  x_G_3_0_m2: CM8 port map (
      D0 => N_7980,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2478,
      D2 => NN_2,
      D3 => NN_2,
      S00 => N_7979,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(57));
  x_G_7_0_m2: CM8 port map (
      D0 => N_7983,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2479,
      D2 => NN_2,
      D3 => NN_2,
      S00 => N_7979,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(56));
  x_G_11_0_m2: CM8 port map (
      D0 => N_7984,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2534,
      D2 => NN_2,
      D3 => NN_2,
      S00 => N_7979,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(1));
  x_I_217: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => rst,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => RST_I);
  x_I_218: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => HOLDN_I);
  x_I_218_0: BUFF port map (
      A => HOLDN_I_0_1,
      Y => HOLDN_I_0);
  x_I_218_0_0: BUFF port map (
      A => HOLDN_I_0_1,
      Y => HOLDN_I_0_0);
  x_I_218_0_1: BUFF port map (
      A => HOLDN_I,
      Y => HOLDN_I_0_1);
  x_I_218_1: BUFF port map (
      A => HOLDN_I_0_1,
      Y => HOLDN_I_1);
  x_I_218_1_0: BUFF port map (
      A => HOLDN_I_0_1,
      Y => HOLDN_I_1_0);
  x_I_218_2: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_2);
  x_I_218_3: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_3);
  x_I_218_4: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_4);
  x_I_218_5: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_5);
  x_I_218_6: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_6);
  x_I_218_7: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_7);
  x_I_218_8: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_8);
  x_I_218_9: BUFF port map (
      A => HOLDN_I_1_0,
      Y => HOLDN_I_9);
  x_I_218_10: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_10);
  x_I_218_11: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_11);
  x_I_218_12: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_12);
  x_I_218_13: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_13);
  x_I_218_14: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_14);
  x_I_218_15: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_15);
  x_I_218_16: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_16);
  x_I_218_17: BUFF port map (
      A => HOLDN_I_0_0,
      Y => HOLDN_I_17);
  NN_3 <= '1';
  x_VCC_Z9647: VCC port map (
      Y => NN_4);
  x_cpi_d_inst_0_31_0x: BUFF port map (
      A => cpi_d_inst(11),
      Y => CPI_D_INST_0(11));
  x_cpi_d_inst_0_0_31_0x: BUFF port map (
      A => cpi_d_inst(9),
      Y => CPI_D_INST_0(9));
  x_cpi_dbg_addr_0_4_0x: BUFF port map (
      A => CPI_DBG_ADDR_0_0(0),
      Y => CPI_DBG_ADDR_0(0));
  x_cpi_dbg_addr_0_0_4_0x: BUFF port map (
      A => cpi_dbg_addr(0),
      Y => CPI_DBG_ADDR_0_0(0));
  x_cpi_dbg_addr_1_4_0x: BUFF port map (
      A => CPI_DBG_ADDR_0_0(0),
      Y => CPI_DBG_ADDR_1(0));
  x_cpi_dbg_addr_2_4_0x: BUFF port map (
      A => CPI_DBG_ADDR_0_0(0),
      Y => CPI_DBG_ADDR_2(0));
  x_cpi_dbg_enable_0: BUFF port map (
      A => cpi_dbg_enable,
      Y => CPI_DBG_ENABLE_0);
  x_cpi_dbg_fsr_0: BUFF port map (
      A => CPI_DBG_FSR_0_0,
      Y => CPI_DBG_FSR_0);
  x_cpi_dbg_fsr_0_0: BUFF port map (
      A => cpi_dbg_fsr,
      Y => CPI_DBG_FSR_0_0);
  x_cpi_dbg_fsr_1: BUFF port map (
      A => CPI_DBG_FSR_0_0,
      Y => CPI_DBG_FSR_1);
  x_cpi_dbg_fsr_2: BUFF port map (
      A => CPI_DBG_FSR_0_0,
      Y => CPI_DBG_FSR_2);
  x_grlfpc2_0_G_167: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_WREN22,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_WREN2_2_SQMUXA_0,
      S01 => cpi_x_inst(20),
      S10 => GRLFPC2_0_WREN1_0_SQMUXA_3,
      S11 => GRLFPC2_0_WREN1_0_SQMUXA_2,
      Y => GRLFPC2_0_N_552);
  x_grlfpc2_0_I_346: AND2B port map (
      A => GRLFPC2_0_R_I_EXEC,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_N_1059);
  x_grlfpc2_0_I_349: CM8 port map (
      D0 => GRLFPC2_0_R_X_SEQERR,
      D1 => GRLFPC2_0_I_349_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1058);
  x_grlfpc2_0_I_349_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_I_EXEC,
      Y => GRLFPC2_0_I_349_CM8I);
  x_grlfpc2_0_I_352: CM8 port map (
      D0 => GRLFPC2_0_I_352_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1,
      S01 => GRLFPC2_0_COMB_CCWR4_1,
      S10 => GRLFPC2_0_COMB_WRRES4,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1063);
  x_grlfpc2_0_I_352_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_COMB_UN3_HOLDN_0,
      S00 => GRLFPC2_0_R_A_MOV,
      S01 => GRLFPC2_0_R_A_FPOP_0,
      S10 => GRLFPC2_0_R_I_EXEC,
      S11 => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_I_352_1);
  x_grlfpc2_0_I_352_2: AND3B port map (
      A => GRLFPC2_0_N_1058,
      B => RST_I,
      C => GRLFPC2_0_I_352_1,
      Y => GRLFPC2_0_I_352_2);
  x_grlfpc2_0_I_352_4: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_COMB_UN1_MEXC,
      S00 => GRLFPC2_0_I_352_2,
      S01 => GRLFPC2_0_ANNULRES_1_SQMUXA_2,
      S10 => GRLFPC2_0_R_I_V,
      S11 => NN_2,
      Y => GRLFPC2_0_I_352_4);
  x_grlfpc2_0_I_361: CM8 port map (
      D0 => GRLFPC2_0_R_I_RDD,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_X_RDD,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_MOV,
      S01 => GRLFPC2_0_COMB_V_E_FPOP_1,
      S10 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1080);
  x_grlfpc2_0_I_378: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_N_1127,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
      S01 => cpi_d_inst(0),
      S10 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
      S11 => GRLFPC2_0_I_378_CM8I,
      Y => GRLFPC2_0_N_1093);
  x_grlfpc2_0_I_378_cm8i: CM8INV port map (
      A => cpi_d_inst(31),
      Y => GRLFPC2_0_I_378_CM8I);
  x_grlfpc2_0_I_382_n: OR2B port map (
      A => cpi_d_inst(14),
      B => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
      Y => GRLFPC2_0_N_1109_N);
  x_grlfpc2_0_I_388: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_N_1109_N,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_FPDECODE_MOV12,
      S01 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
      S10 => GRLFPC2_0_COMB_FPDECODE_MOV12,
      S11 => GRLFPC2_0_I_388_CM8I,
      Y => GRLFPC2_0_N_1108);
  x_grlfpc2_0_I_388_cm8i: CM8INV port map (
      A => GRLFPC2_0_RS1D_CNST,
      Y => GRLFPC2_0_I_388_CM8I);
  x_grlfpc2_0_I_391: CM8 port map (
      D0 => NN_2,
      D1 => cpi_d_inst(25),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_N_1105,
      S01 => cpi_d_inst(31),
      S10 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      S11 => GRLFPC2_0_N_335,
      Y => GRLFPC2_0_N_1104);
  x_grlfpc2_0_I_394: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_RS1V10,
      D2 => NN_2,
      D3 => GRLFPC2_0_RS1V10,
      S00 => cpi_d_inst(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_N_1108,
      S11 => GRLFPC2_0_N_353_1,
      Y => GRLFPC2_0_N_1105);
  x_grlfpc2_0_I_402: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      D2 => cpi_d_inst(0),
      D3 => NN_4,
      S00 => GRLFPC2_0_N_1127,
      S01 => NN_4,
      S10 => GRLFPC2_0_RS2_0_SQMUXA,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1123);
  x_grlfpc2_0_I_406: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
      D2 => GRLFPC2_0_COMB_FPDECODE_MOV11,
      D3 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
      S00 => GRLFPC2_0_COMB_FPDECODE_MOV12,
      S01 => NN_4,
      S10 => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_1,
      S11 => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210,
      Y => GRLFPC2_0_N_1127);
  x_grlfpc2_0_I_416: AND3A port map (
      A => GRLFPC2_0_RS1D_CNST,
      B => cpi_d_inst(25),
      C => cpi_d_inst(30),
      Y => GRLFPC2_0_N_1133);
  x_grlfpc2_0_I_422: CM8 port map (
      D0 => NN_4,
      D1 => cpi_d_inst(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_I_423_0,
      S01 => GRLFPC2_0_N_816,
      S10 => GRLFPC2_0_N_1133,
      S11 => GRLFPC2_0_I_422_CM8I,
      Y => GRLFPC2_0_N_1132);
  x_grlfpc2_0_I_422_1_n: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_I_422_1_N_CM8I,
      D2 => NN_2,
      D3 => GRLFPC2_0_RS1V10,
      S00 => cpi_d_inst(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1132_1_N);
  x_grlfpc2_0_I_422_1_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_N_353_1,
      Y => GRLFPC2_0_I_422_1_N_CM8I);
  x_grlfpc2_0_I_422_cm8i: CM8INV port map (
      A => GRLFPC2_0_N_1132_1_N,
      Y => GRLFPC2_0_I_422_CM8I);
  x_grlfpc2_0_I_423_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_FPDECODE_MOV12,
      S01 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
      S10 => GRLFPC2_0_COMB_FPDECODE_MOV12,
      S11 => GRLFPC2_0_I_423_0_CM8I,
      Y => GRLFPC2_0_I_423_0);
  x_grlfpc2_0_I_423_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_RS1D_CNST,
      Y => GRLFPC2_0_I_423_0_CM8I);
  x_grlfpc2_0_annulres_0_sqmuxa_3_1: AND4B port map (
      A => GRLFPC2_0_R_M_FPOP,
      B => GRLFPC2_0_R_E_FPOP,
      C => GRLFPC2_0_R_A_FPOP_0,
      D => GRLFPC2_0_COMB_UN3_HOLDN_0,
      Y => GRLFPC2_0_ANNULRES_0_SQMUXA_3_1);
  x_grlfpc2_0_annulres_0_sqmuxa_4_1: AND2A port map (
      A => GRLFPC2_0_R_I_EXEC,
      B => GRLFPC2_0_R_X_FPOP,
      Y => GRLFPC2_0_ANNULRES_0_SQMUXA_4_1);
  x_grlfpc2_0_annulres_1_sqmuxa_2: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_ANNULRES_0_SQMUXA_3_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_N_1059,
      S11 => NN_2,
      Y => GRLFPC2_0_ANNULRES_1_SQMUXA_2);
  x_grlfpc2_0_annulres_1_sqmuxa_2_tz_0: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0_CM8I,
      D3 => GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0_CM8I,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_2,
      S01 => GRLFPC2_0_R_E_FPOP,
      S10 => GRLFPC2_0_R_M_FPOP,
      S11 => NN_2,
      Y => GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0);
  x_grlfpc2_0_annulres_1_sqmuxa_2_tz_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1,
      Y => GRLFPC2_0_ANNULRES_1_SQMUXA_2_TZ_0_CM8I);
  x_grlfpc2_0_comb_annulfpu_1_0: CM8 port map (
      D0 => GRLFPC2_0_R_X_SEQERR,
      D1 => GRLFPC2_0_R_X_FPOP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_849);
  x_grlfpc2_0_comb_annulfpu_1_u: CM8 port map (
      D0 => GRLFPC2_0_COMB_ANNULFPU_1_U_0,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_1,
      S01 => GRLFPC2_0_R_M_FPOP,
      S10 => GRLFPC2_0_N_849,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_ANNULFPU_1);
  x_grlfpc2_0_comb_annulfpu_1_u_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_R_A_FPOP,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_2,
      S01 => GRLFPC2_0_R_E_FPOP,
      S10 => GRLFPC2_0_COMB_UN3_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_ANNULFPU_1_U_0);
  x_grlfpc2_0_comb_annulres_1: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_UN1_FPCI_3_1,
      D2 => NN_4,
      D3 => GRLFPC2_0_ANNULRES_0_SQMUXA_4_1,
      S00 => GRLFPC2_0_ANNULRES_1_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_ANNULRES_1);
  x_grlfpc2_0_comb_ccwr4_1: AND2A port map (
      A => GRLFPC2_0_COMB_V_STATE_7(0),
      B => GRLFPC2_0_COMB_CCWR4_1_0,
      Y => GRLFPC2_0_COMB_CCWR4_1);
  x_grlfpc2_0_comb_ccwr4_1_0: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_V_I_V6,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_R_I_V,
      S01 => GRLFPC2_0_COMB_V_I_EXEC_4,
      S10 => GRLFPC2_0_COMB_CCWR4_1_0_CM8I,
      S11 => GRLFPC2_0_UN1_FPCI_2_N,
      Y => GRLFPC2_0_COMB_CCWR4_1_0);
  x_grlfpc2_0_comb_ccwr4_1_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_STATE(1),
      Y => GRLFPC2_0_COMB_CCWR4_1_0_CM8I);
  x_grlfpc2_0_comb_dbgdata_5_0x: CM8 port map (
      D0 => rfo1_data1(0),
      D1 => GRLFPC2_0_R_FSR_CEXC(0),
      D2 => rfo2_data1(0),
      D3 => GRLFPC2_0_R_FSR_CEXC(0),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(0));
  x_grlfpc2_0_comb_dbgdata_5_1x: CM8 port map (
      D0 => rfo1_data1(1),
      D1 => GRLFPC2_0_R_FSR_CEXC(1),
      D2 => rfo2_data1(1),
      D3 => GRLFPC2_0_R_FSR_CEXC(1),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(1));
  x_grlfpc2_0_comb_dbgdata_5_2x: CM8 port map (
      D0 => rfo1_data1(2),
      D1 => GRLFPC2_0_R_FSR_CEXC(2),
      D2 => rfo2_data1(2),
      D3 => GRLFPC2_0_R_FSR_CEXC(2),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(2));
  x_grlfpc2_0_comb_dbgdata_5_3x: CM8 port map (
      D0 => rfo1_data1(3),
      D1 => GRLFPC2_0_R_FSR_CEXC(3),
      D2 => rfo2_data1(3),
      D3 => GRLFPC2_0_R_FSR_CEXC(3),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(3));
  x_grlfpc2_0_comb_dbgdata_5_4x: CM8 port map (
      D0 => rfo1_data1(4),
      D1 => GRLFPC2_0_R_FSR_CEXC(4),
      D2 => rfo2_data1(4),
      D3 => GRLFPC2_0_R_FSR_CEXC(4),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(4));
  x_grlfpc2_0_comb_dbgdata_5_5x: CM8 port map (
      D0 => rfo1_data1(5),
      D1 => GRLFPC2_0_R_FSR_AEXC(0),
      D2 => rfo2_data1(5),
      D3 => GRLFPC2_0_R_FSR_AEXC(0),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(5));
  x_grlfpc2_0_comb_dbgdata_5_6x: CM8 port map (
      D0 => rfo1_data1(6),
      D1 => GRLFPC2_0_R_FSR_AEXC(1),
      D2 => rfo2_data1(6),
      D3 => GRLFPC2_0_R_FSR_AEXC(1),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(6));
  x_grlfpc2_0_comb_dbgdata_5_7x: CM8 port map (
      D0 => rfo1_data1(7),
      D1 => GRLFPC2_0_R_FSR_AEXC(2),
      D2 => rfo2_data1(7),
      D3 => GRLFPC2_0_R_FSR_AEXC(2),
      S00 => CPI_DBG_FSR_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(7));
  x_grlfpc2_0_comb_dbgdata_5_8x: CM8 port map (
      D0 => rfo1_data1(8),
      D1 => GRLFPC2_0_R_FSR_AEXC(3),
      D2 => rfo2_data1(8),
      D3 => GRLFPC2_0_R_FSR_AEXC(3),
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(8));
  x_grlfpc2_0_comb_dbgdata_5_9x: CM8 port map (
      D0 => rfo1_data1(9),
      D1 => GRLFPC2_0_R_FSR_AEXC(4),
      D2 => rfo2_data1(9),
      D3 => GRLFPC2_0_R_FSR_AEXC(4),
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(9));
  x_grlfpc2_0_comb_dbgdata_5_10x: CM8 port map (
      D0 => rfo1_data1(10),
      D1 => CPO_CC_0_INT_2,
      D2 => rfo2_data1(10),
      D3 => CPO_CC_0_INT_2,
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(10));
  x_grlfpc2_0_comb_dbgdata_5_11x: CM8 port map (
      D0 => rfo1_data1(11),
      D1 => CPO_CC_1_INT_3,
      D2 => rfo2_data1(11),
      D3 => CPO_CC_1_INT_3,
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(11));
  x_grlfpc2_0_comb_dbgdata_5_12x: CM8 port map (
      D0 => rfo1_data1(12),
      D1 => NN_2,
      D2 => rfo2_data1(12),
      D3 => NN_2,
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(12));
  x_grlfpc2_0_comb_dbgdata_5_13x: CM8 port map (
      D0 => rfo1_data1(13),
      D1 => GRLFPC2_0_COMB_QNE2,
      D2 => rfo2_data1(13),
      D3 => GRLFPC2_0_COMB_QNE2,
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(13));
  x_grlfpc2_0_comb_dbgdata_5_14x: CM8 port map (
      D0 => rfo1_data1(14),
      D1 => GRLFPC2_0_R_FSR_FTT(0),
      D2 => rfo2_data1(14),
      D3 => GRLFPC2_0_R_FSR_FTT(0),
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(14));
  x_grlfpc2_0_comb_dbgdata_5_15x: CM8 port map (
      D0 => rfo1_data1(15),
      D1 => NN_2,
      D2 => rfo2_data1(15),
      D3 => NN_2,
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(15));
  x_grlfpc2_0_comb_dbgdata_5_16x: CM8 port map (
      D0 => rfo1_data1(16),
      D1 => GRLFPC2_0_R_FSR_FTT(2),
      D2 => rfo2_data1(16),
      D3 => GRLFPC2_0_R_FSR_FTT(2),
      S00 => CPI_DBG_FSR_1,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(16));
  x_grlfpc2_0_comb_dbgdata_5_17x: CM8 port map (
      D0 => rfo1_data1(17),
      D1 => NN_4,
      D2 => rfo2_data1(17),
      D3 => NN_4,
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_1(0),
      S11 => NN_2,
      Y => cpo_dbg_data(17));
  x_grlfpc2_0_comb_dbgdata_5_18x: CM8 port map (
      D0 => rfo1_data1(18),
      D1 => NN_4,
      D2 => rfo2_data1(18),
      D3 => NN_4,
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(18));
  x_grlfpc2_0_comb_dbgdata_5_19x: CM8 port map (
      D0 => rfo1_data1(19),
      D1 => NN_2,
      D2 => rfo2_data1(19),
      D3 => NN_2,
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(19));
  x_grlfpc2_0_comb_dbgdata_5_20x: CM8 port map (
      D0 => rfo1_data1(20),
      D1 => NN_2,
      D2 => rfo2_data1(20),
      D3 => NN_2,
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(20));
  x_grlfpc2_0_comb_dbgdata_5_21x: CM8 port map (
      D0 => rfo1_data1(21),
      D1 => NN_2,
      D2 => rfo2_data1(21),
      D3 => NN_2,
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(21));
  x_grlfpc2_0_comb_dbgdata_5_22x: CM8 port map (
      D0 => rfo1_data1(22),
      D1 => GRLFPC2_0_R_FSR_NONSTD,
      D2 => rfo2_data1(22),
      D3 => GRLFPC2_0_R_FSR_NONSTD,
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(22));
  x_grlfpc2_0_comb_dbgdata_5_23x: CM8 port map (
      D0 => rfo1_data1(23),
      D1 => GRLFPC2_0_R_FSR_TEM(0),
      D2 => rfo2_data1(23),
      D3 => GRLFPC2_0_R_FSR_TEM(0),
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(23));
  x_grlfpc2_0_comb_dbgdata_5_24x: CM8 port map (
      D0 => rfo1_data1(24),
      D1 => GRLFPC2_0_R_FSR_TEM(1),
      D2 => rfo2_data1(24),
      D3 => GRLFPC2_0_R_FSR_TEM(1),
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(24));
  x_grlfpc2_0_comb_dbgdata_5_25x: CM8 port map (
      D0 => rfo1_data1(25),
      D1 => GRLFPC2_0_R_FSR_TEM(2),
      D2 => rfo2_data1(25),
      D3 => GRLFPC2_0_R_FSR_TEM(2),
      S00 => CPI_DBG_FSR_2,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(25));
  x_grlfpc2_0_comb_dbgdata_5_26x: CM8 port map (
      D0 => rfo1_data1(26),
      D1 => GRLFPC2_0_R_FSR_TEM(3),
      D2 => rfo2_data1(26),
      D3 => GRLFPC2_0_R_FSR_TEM(3),
      S00 => CPI_DBG_FSR_0_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_2(0),
      S11 => NN_2,
      Y => cpo_dbg_data(26));
  x_grlfpc2_0_comb_dbgdata_5_27x: CM8 port map (
      D0 => rfo1_data1(27),
      D1 => GRLFPC2_0_R_FSR_TEM(4),
      D2 => rfo2_data1(27),
      D3 => GRLFPC2_0_R_FSR_TEM(4),
      S00 => CPI_DBG_FSR_0_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(27));
  x_grlfpc2_0_comb_dbgdata_5_28x: CM8 port map (
      D0 => rfo1_data1(28),
      D1 => NN_2,
      D2 => rfo2_data1(28),
      D3 => NN_2,
      S00 => CPI_DBG_FSR_0_0,
      S01 => NN_4,
      S10 => CPI_DBG_ADDR_0_0(0),
      S11 => NN_2,
      Y => cpo_dbg_data(28));
  x_grlfpc2_0_comb_dbgdata_5_29x: CM8 port map (
      D0 => rfo1_data1(29),
      D1 => NN_2,
      D2 => rfo2_data1(29),
      D3 => NN_2,
      S00 => cpi_dbg_fsr,
      S01 => NN_4,
      S10 => cpi_dbg_addr(0),
      S11 => NN_2,
      Y => cpo_dbg_data(29));
  x_grlfpc2_0_comb_dbgdata_5_30x: CM8 port map (
      D0 => rfo1_data1(30),
      D1 => GRLFPC2_0_R_FSR_RD(0),
      D2 => rfo2_data1(30),
      D3 => GRLFPC2_0_R_FSR_RD(0),
      S00 => cpi_dbg_fsr,
      S01 => NN_4,
      S10 => cpi_dbg_addr(0),
      S11 => NN_2,
      Y => cpo_dbg_data(30));
  x_grlfpc2_0_comb_dbgdata_5_31x: CM8 port map (
      D0 => rfo1_data1(31),
      D1 => GRLFPC2_0_R_FSR_RD(1),
      D2 => rfo2_data1(31),
      D3 => GRLFPC2_0_R_FSR_RD(1),
      S00 => cpi_dbg_fsr,
      S01 => NN_4,
      S10 => cpi_dbg_addr(0),
      S11 => NN_2,
      Y => cpo_dbg_data(31));
  x_grlfpc2_0_comb_fpdecode_afq3: AND3 port map (
      A => GRLFPC2_0_COMB_FPDECODE_AFQ3_1,
      B => GRLFPC2_0_COMB_RDD_1_1,
      C => GRLFPC2_0_N_17_1,
      Y => GRLFPC2_0_COMB_FPDECODE_AFQ3);
  x_grlfpc2_0_comb_fpdecode_afq3_1: AND2 port map (
      A => cpi_d_inst(21),
      B => cpi_d_inst(20),
      Y => GRLFPC2_0_COMB_FPDECODE_AFQ3_1);
  x_grlfpc2_0_comb_fpdecode_afq6_n: CM8 port map (
      D0 => NN_4,
      D1 => cpi_d_inst(23),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_FPDECODE_AFQ6_N_CM8I,
      S01 => GRLFPC2_0_COMB_RDD_1_1,
      S10 => GRLFPC2_0_COMB_FPDECODE_ST_1,
      S11 => cpi_d_inst(20),
      Y => GRLFPC2_0_COMB_FPDECODE_AFQ6_N);
  x_grlfpc2_0_comb_fpdecode_afq6_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_N_17_1,
      Y => GRLFPC2_0_COMB_FPDECODE_AFQ6_N_CM8I);
  x_grlfpc2_0_comb_fpdecode_afq12: AND2A port map (
      A => cpi_d_inst(30),
      B => cpi_d_inst(31),
      Y => GRLFPC2_0_COMB_FPDECODE_AFQ12);
  x_grlfpc2_0_comb_fpdecode_afq13: AND2 port map (
      A => cpi_d_inst(31),
      B => cpi_d_inst(30),
      Y => GRLFPC2_0_COMB_FPDECODE_AFQ13);
  x_grlfpc2_0_comb_fpdecode_mov2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_MOV2_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_FPDECODE_MOV2_CM8I,
      S01 => cpi_d_inst(12),
      S10 => CPI_D_INST_0(9),
      S11 => cpi_d_inst(6),
      Y => GRLFPC2_0_COMB_FPDECODE_MOV2);
  x_grlfpc2_0_comb_fpdecode_mov2_0: AND2 port map (
      A => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_4,
      B => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV2_0);
  x_grlfpc2_0_comb_fpdecode_mov2_cm8i: CM8INV port map (
      A => cpi_d_inst(10),
      Y => GRLFPC2_0_COMB_FPDECODE_MOV2_CM8I);
  x_grlfpc2_0_comb_fpdecode_mov4_2: AND4C port map (
      A => cpi_d_inst(5),
      B => cpi_d_inst(13),
      C => CPI_D_INST_0(9),
      D => cpi_d_inst(6),
      Y => GRLFPC2_0_COMB_FPDECODE_MOV4_2);
  x_grlfpc2_0_comb_fpdecode_mov5: AND3A port map (
      A => CPI_D_INST_0(9),
      B => GRLFPC2_0_COMB_FPDECODE_MOV5_1,
      C => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV5);
  x_grlfpc2_0_comb_fpdecode_mov5_1: AND3A port map (
      A => cpi_d_inst(5),
      B => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
      C => cpi_d_inst(6),
      Y => GRLFPC2_0_COMB_FPDECODE_MOV5_1);
  x_grlfpc2_0_comb_fpdecode_mov6: AND4A port map (
      A => CPI_D_INST_0(9),
      B => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_3,
      C => GRLFPC2_0_COMB_FPDECODE_MOV4_3,
      D => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV6);
  x_grlfpc2_0_comb_fpdecode_mov6_2: AND3B port map (
      A => cpi_d_inst(12),
      B => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2,
      C => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_4,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV4_3);
  x_grlfpc2_0_comb_fpdecode_mov7: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1,
      D1 => NN_4,
      D2 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1,
      D3 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1,
      S00 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_4,
      S01 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_3,
      S10 => GRLFPC2_0_COMB_FPDECODE_MOV7_CM8I,
      S11 => CPI_D_INST_0(11),
      Y => GRLFPC2_0_COMB_FPDECODE_MOV7);
  x_grlfpc2_0_comb_fpdecode_mov7_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_5,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV7_CM8I);
  x_grlfpc2_0_comb_fpdecode_mov11: AND4B port map (
      A => GRLFPC2_0_COMB_FPDECODE_ST_1,
      B => cpi_d_inst(19),
      C => GRLFPC2_0_COMB_RDD_1_1,
      D => GRLFPC2_0_N_16_1,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV11);
  x_grlfpc2_0_comb_fpdecode_mov12: AND2 port map (
      A => cpi_d_inst(19),
      B => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
      Y => GRLFPC2_0_COMB_FPDECODE_MOV12);
  x_grlfpc2_0_comb_fpdecode_rs2d5: AND2 port map (
      A => GRLFPC2_0_COMB_FPDECODE_RS2D5_0,
      B => GRLFPC2_0_COMB_FPDECODE_MOV5_1,
      Y => GRLFPC2_0_COMB_FPDECODE_RS2D5);
  x_grlfpc2_0_comb_fpdecode_rs2d5_0: AND3A port map (
      A => cpi_d_inst(8),
      B => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2,
      C => CPI_D_INST_0(9),
      Y => GRLFPC2_0_COMB_FPDECODE_RS2D5_0);
  x_grlfpc2_0_comb_fpdecode_rs2d5_1: AND2A port map (
      A => cpi_d_inst(13),
      B => CPI_D_INST_0(11),
      Y => GRLFPC2_0_COMB_FPDECODE_RS2D5_1);
  x_grlfpc2_0_comb_fpdecode_st_0_a2: AND2 port map (
      A => GRLFPC2_0_COMB_FPDECODE_ST_1,
      B => GRLFPC2_0_COMB_V_A_AFQ_1_1_0,
      Y => GRLFPC2_0_COMB_FPDECODE_ST);
  x_grlfpc2_0_comb_fpdecode_st_0_a2_1: AND2A port map (
      A => cpi_d_inst(23),
      B => cpi_d_inst(21),
      Y => GRLFPC2_0_COMB_FPDECODE_ST_1);
  x_grlfpc2_0_comb_fpdecode_un1_fpci_1: AND4B port map (
      A => CPI_D_INST_0(11),
      B => cpi_d_inst(8),
      C => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_5,
      D => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_3,
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1);
  x_grlfpc2_0_comb_fpdecode_un1_fpci_1_2: AND3B port map (
      A => CPI_D_INST_0(9),
      B => cpi_d_inst(13),
      C => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2,
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_5);
  x_grlfpc2_0_comb_fpdecode_un1_fpci_2: AND2B port map (
      A => cpi_d_inst(10),
      B => cpi_d_inst(12),
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2);
  x_grlfpc2_0_comb_fpdecode_un1_fpci_3: AND2A port map (
      A => cpi_d_inst(6),
      B => cpi_d_inst(5),
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_3);
  x_grlfpc2_0_comb_fpdecode_un1_fpci_4: AND2A port map (
      A => cpi_d_inst(7),
      B => cpi_d_inst(8),
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_4);
  x_grlfpc2_0_comb_fpdecode_un1_wren210: AND2A port map (
      A => cpi_d_inst(7),
      B => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0,
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210);
  x_grlfpc2_0_comb_fpdecode_un1_wren210_1_0: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_MOV5_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0_CM8I,
      S01 => CPI_D_INST_0(9),
      S10 => cpi_d_inst(8),
      S11 => cpi_d_inst(10),
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0);
  x_grlfpc2_0_comb_fpdecode_un1_wren210_1_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_FPDECODE_RS2D5_0,
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0_CM8I);
  x_grlfpc2_0_comb_fpdecode_un1_wren210_1_1_0: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_MOV4_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => CPI_D_INST_0(11),
      S01 => cpi_d_inst(7),
      S10 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2,
      S11 => cpi_d_inst(10),
      Y => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_1_0);
  x_grlfpc2_0_comb_fpdecode_un3_op: AND3 port map (
      A => cpi_d_inst(23),
      B => GRLFPC2_0_COMB_RDD_1_1,
      C => GRLFPC2_0_N_16_1,
      Y => GRLFPC2_0_COMB_FPDECODE_UN3_OP);
  x_grlfpc2_0_comb_fpop_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN4_LOCK,
      B => GRLFPC2_0_RS2_0_SQMUXA,
      Y => GRLFPC2_0_COMB_FPOP_1);
  x_grlfpc2_0_comb_isfpop2_1: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(19),
      D1 => cpi_x_inst(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1_CM8I,
      S01 => GRLFPC2_0_R_X_FPOP,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_ISFPOP2_1);
  x_grlfpc2_0_comb_isfpop2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_I_EXEC,
      Y => GRLFPC2_0_COMB_ISFPOP2_1_CM8I);
  x_grlfpc2_0_comb_lock_1: AND4C port map (
      A => GRLFPC2_0_N_331,
      B => cpi_d_trap,
      C => cpi_d_annul,
      D => GRLFPC2_0_COMB_LOCK_1_0,
      Y => cpo_ldlock);
  x_grlfpc2_0_comb_lock_1_0: AND2B port map (
      A => GRLFPC2_0_R_STATE(0),
      B => GRLFPC2_0_R_STATE(1),
      Y => GRLFPC2_0_COMB_LOCK_1_0);
  x_grlfpc2_0_comb_lockgen_depcheck: OR4 port map (
      A => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK_1,
      B => GRLFPC2_0_R_X_FPOP,
      C => GRLFPC2_0_R_A_FPOP,
      D => GRLFPC2_0_R_E_FPOP,
      Y => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK);
  x_grlfpc2_0_comb_lockgen_depcheck_1: OR2 port map (
      A => GRLFPC2_0_R_M_FPOP,
      B => GRLFPC2_0_R_I_EXEC,
      Y => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK_1);
  x_grlfpc2_0_comb_lockgen_locki_i: CM8 port map (
      D0 => GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_CM8I,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_LOCKGEN_UN6_DEPCHECK,
      S01 => GRLFPC2_0_COMB_LOCKGEN_UN8_DEPCHECK,
      S10 => GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_1,
      S11 => NN_2,
      Y => GRLFPC2_0_N_331);
  x_grlfpc2_0_comb_lockgen_locki_i_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => cpi_d_cnt(0),
      D3 => NN_4,
      S00 => cpi_d_cnt(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_SEQERR_UN7_OP,
      S11 => GRLFPC2_0_COMB_FPDECODE_ST,
      Y => GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_1);
  x_grlfpc2_0_comb_lockgen_locki_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK,
      Y => GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_CM8I);
  x_grlfpc2_0_comb_lockgen_un6_depcheck: OR2 port map (
      A => GRLFPC2_0_RS2_0_SQMUXA,
      B => GRLFPC2_0_COMB_FPDECODE_ST,
      Y => GRLFPC2_0_COMB_LOCKGEN_UN6_DEPCHECK);
  x_grlfpc2_0_comb_lockgen_un8_depcheck: OR4 port map (
      A => GRLFPC2_0_R_X_LD_0,
      B => GRLFPC2_0_R_M_LD,
      C => GRLFPC2_0_R_E_LD,
      D => GRLFPC2_0_R_A_LD,
      Y => GRLFPC2_0_COMB_LOCKGEN_UN8_DEPCHECK);
  x_grlfpc2_0_comb_mexc_1_1x: AND2 port map (
      A => GRLFPC2_0_R_I_EXC(1),
      B => GRLFPC2_0_R_FSR_TEM(1),
      Y => GRLFPC2_0_COMB_MEXC_1(1));
  x_grlfpc2_0_comb_mexc_1_2x: AND2 port map (
      A => GRLFPC2_0_R_I_EXC(2),
      B => GRLFPC2_0_R_FSR_TEM(2),
      Y => GRLFPC2_0_COMB_MEXC_1(2));
  x_grlfpc2_0_comb_pexc9: AND2A port map (
      A => GRLFPC2_0_R_STATE(1),
      B => GRLFPC2_0_R_STATE(0),
      Y => CPO_EXC_INT_1);
  x_grlfpc2_0_comb_qne2: AND2A port map (
      A => GRLFPC2_0_R_STATE(0),
      B => GRLFPC2_0_R_STATE(1),
      Y => GRLFPC2_0_COMB_QNE2);
  x_grlfpc2_0_comb_rdd_3: CM8 port map (
      D0 => GRLFPC2_0_R_I_RDD,
      D1 => GRLFPC2_0_R_I_RDD,
      D2 => GRLFPC2_0_R_I_RDD,
      D3 => GRLFPC2_0_R_X_RDD,
      S00 => GRLFPC2_0_ANNULRES_0_SQMUXA_4_1,
      S01 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S10 => GRLFPC2_0_R_I_V,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RDD_3);
  x_grlfpc2_0_comb_rdd_3_0: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_0);
  x_grlfpc2_0_comb_rdd_3_0_0: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3,
      Y => GRLFPC2_0_COMB_RDD_3_0_0);
  x_grlfpc2_0_comb_rdd_3_1: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_1);
  x_grlfpc2_0_comb_rdd_3_2: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_2);
  x_grlfpc2_0_comb_rdd_3_3: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_3);
  x_grlfpc2_0_comb_rdd_3_4: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_4);
  x_grlfpc2_0_comb_rdd_3_5: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_5);
  x_grlfpc2_0_comb_rdd_3_6: BUFF port map (
      A => GRLFPC2_0_COMB_RDD_3_0_0,
      Y => GRLFPC2_0_COMB_RDD_3_6);
  x_grlfpc2_0_comb_rs1_1_0x: CM8 port map (
      D0 => GRLFPC2_0_N_816,
      D1 => NN_2,
      D2 => GRLFPC2_0_N_816,
      D3 => cpi_d_inst(25),
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_RS1V_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS1_1(0));
  x_grlfpc2_0_comb_rs1_1_1x: CM8 port map (
      D0 => GRLFPC2_0_N_817,
      D1 => NN_2,
      D2 => GRLFPC2_0_N_817,
      D3 => cpi_d_inst(26),
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_RS1V_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS1_1(1));
  x_grlfpc2_0_comb_rs1_1_2x: CM8 port map (
      D0 => GRLFPC2_0_N_818,
      D1 => NN_2,
      D2 => GRLFPC2_0_N_818,
      D3 => cpi_d_inst(27),
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_RS1V_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS1_1(2));
  x_grlfpc2_0_comb_rs1_1_3x: CM8 port map (
      D0 => GRLFPC2_0_N_819,
      D1 => NN_2,
      D2 => GRLFPC2_0_N_819,
      D3 => cpi_d_inst(28),
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_RS1V_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS1_1(3));
  x_grlfpc2_0_comb_rs1_1_4x: CM8 port map (
      D0 => GRLFPC2_0_N_820,
      D1 => NN_2,
      D2 => GRLFPC2_0_N_820,
      D3 => cpi_d_inst(29),
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_RS1V_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS1_1(4));
  x_grlfpc2_0_comb_rs1_1_0_0x: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(0),
      D1 => cpi_d_inst(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_816);
  x_grlfpc2_0_comb_rs1_1_0_1x: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(1),
      D1 => cpi_d_inst(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_817);
  x_grlfpc2_0_comb_rs1_1_0_2x: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(2),
      D1 => cpi_d_inst(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_818);
  x_grlfpc2_0_comb_rs1_1_0_3x: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(3),
      D1 => cpi_d_inst(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_819);
  x_grlfpc2_0_comb_rs1_1_0_4x: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(4),
      D1 => cpi_d_inst(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_820);
  x_grlfpc2_0_comb_rs1d_1_u: CM8 port map (
      D0 => GRLFPC2_0_RS1D_CNST,
      D1 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_MOV_7_SQMUXA,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS1D_1);
  x_grlfpc2_0_comb_rs1v_1_i_a4_0_1: AND2A port map (
      A => GRLFPC2_0_COMB_FPDECODE_MOV5,
      B => GRLFPC2_0_COMB_RS1V_1_I_A4_0_1_1,
      Y => GRLFPC2_0_N_353_1);
  x_grlfpc2_0_comb_rs1v_1_i_a4_0_1_0: AND2A port map (
      A => GRLFPC2_0_COMB_RSDECODE_UN1_FPCI,
      B => GRLFPC2_0_COMB_FPDECODE_MOV11,
      Y => GRLFPC2_0_COMB_RS1V_1_I_A4_0_1_0);
  x_grlfpc2_0_comb_rs1v_1_i_a4_0_1_1: AND2A port map (
      A => GRLFPC2_0_COMB_FPDECODE_MOV6,
      B => GRLFPC2_0_COMB_RS1V_1_I_A4_0_1_0,
      Y => GRLFPC2_0_COMB_RS1V_1_I_A4_0_1_1);
  x_grlfpc2_0_comb_rs2_1_0x: CM8 port map (
      D0 => cpi_d_inst(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS2(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => HOLDN_I_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_RS2_1(0));
  x_grlfpc2_0_comb_rs2_1_1x: CM8 port map (
      D0 => cpi_d_inst(1),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2_0,
      S01 => NN_4,
      S10 => HOLDN_I_1,
      S11 => NN_2,
      Y => RFI2_RD2ADDR_0_INT_9_INT_22);
  x_grlfpc2_0_comb_rs2_1_2x: CM8 port map (
      D0 => cpi_d_inst(2),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      S01 => NN_4,
      S10 => HOLDN_I_1,
      S11 => NN_2,
      Y => RFI2_RD2ADDR_1_INT_10_INT_23);
  x_grlfpc2_0_comb_rs2_1_3x: CM8 port map (
      D0 => cpi_d_inst(3),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      S01 => NN_4,
      S10 => HOLDN_I_1,
      S11 => NN_2,
      Y => RFI2_RD2ADDR_2_INT_11_INT_24);
  x_grlfpc2_0_comb_rs2_1_4x: CM8 port map (
      D0 => cpi_d_inst(4),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS2(4),
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      S01 => NN_4,
      S10 => HOLDN_I_1,
      S11 => NN_2,
      Y => RFI2_RD2ADDR_3_INT_12_INT_25);
  x_grlfpc2_0_comb_rs2_1_sn_m1: AND2B port map (
      A => HOLDN_I_1,
      B => GRLFPC2_0_RS2_0_SQMUXA,
      Y => GRLFPC2_0_COMB_RS2_1_SN_N_2);
  x_grlfpc2_0_comb_rs2_1_sn_m1_0: AND2B port map (
      A => HOLDN_I_1,
      B => GRLFPC2_0_RS2_0_SQMUXA,
      Y => GRLFPC2_0_COMB_RS2_1_SN_N_2_0);
  x_grlfpc2_0_comb_rs2d_1: AND2 port map (
      A => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      B => GRLFPC2_0_N_1127,
      Y => GRLFPC2_0_COMB_RS2D_1);
  x_grlfpc2_0_comb_rsdecode_un1_fpci: AND4A port map (
      A => cpi_d_inst(9),
      B => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_3,
      C => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_2,
      D => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
      Y => GRLFPC2_0_COMB_RSDECODE_UN1_FPCI);
  x_grlfpc2_0_comb_seqerr_un7_op: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_SEQERR_UN7_OP_CM8I,
      S01 => GRLFPC2_0_COMB_FPDECODE_AFQ6_N,
      S10 => GRLFPC2_0_RS2_0_SQMUXA,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_SEQERR_UN7_OP);
  x_grlfpc2_0_comb_seqerr_un7_op_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_SEQERR_UN11_OP_0,
      Y => GRLFPC2_0_COMB_SEQERR_UN7_OP_CM8I);
  x_grlfpc2_0_comb_seqerr_un11_op_0: AND3A port map (
      A => GRLFPC2_0_COMB_FPDECODE_ST_1,
      B => GRLFPC2_0_N_17_1,
      C => GRLFPC2_0_COMB_RDD_1_1,
      Y => GRLFPC2_0_COMB_SEQERR_UN11_OP_0);
  x_grlfpc2_0_comb_un1_fpci: OR3 port map (
      A => cpi_flush,
      B => cpi_x_annul,
      C => cpi_x_trap,
      Y => GRLFPC2_0_COMB_UN1_FPCI);
  x_grlfpc2_0_comb_un1_fpci_0: OR3 port map (
      A => cpi_flush,
      B => cpi_x_annul,
      C => cpi_x_trap,
      Y => GRLFPC2_0_COMB_UN1_FPCI_0);
  x_grlfpc2_0_comb_un1_fpci_1: OR2 port map (
      A => cpi_m_trap,
      B => cpi_m_annul,
      Y => GRLFPC2_0_COMB_UN1_FPCI_1);
  x_grlfpc2_0_comb_un1_fpci_1_0: OR3 port map (
      A => cpi_flush,
      B => cpi_x_annul,
      C => cpi_x_trap,
      Y => GRLFPC2_0_COMB_UN1_FPCI_1_0);
  x_grlfpc2_0_comb_un1_fpci_2: OR2 port map (
      A => cpi_e_trap,
      B => cpi_e_annul,
      Y => GRLFPC2_0_COMB_UN1_FPCI_2);
  x_grlfpc2_0_comb_un1_fpci_3: AND3 port map (
      A => GRLFPC2_0_R_A_RS1D,
      B => cpi_a_cnt(1),
      C => GRLFPC2_0_R_A_ST,
      Y => GRLFPC2_0_COMB_UN1_FPCI_3);
  x_grlfpc2_0_comb_un1_fpci_4: CM8 port map (
      D0 => GRLFPC2_0_COMB_UN1_FPCI_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_CM8I,
      S01 => GRLFPC2_0_R_A_RS2(0),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4);
  x_grlfpc2_0_comb_un1_fpci_4_0: CM8 port map (
      D0 => GRLFPC2_0_COMB_UN1_FPCI_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0_CM8I,
      S01 => GRLFPC2_0_R_A_RS2(0),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_0);
  x_grlfpc2_0_comb_un1_fpci_4_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_A_RS2D,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_0_CM8I);
  x_grlfpc2_0_comb_un1_fpci_4_1: CM8 port map (
      D0 => GRLFPC2_0_COMB_UN1_FPCI_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1_CM8I,
      S01 => GRLFPC2_0_R_A_RS2(0),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_1);
  x_grlfpc2_0_comb_un1_fpci_4_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_A_RS2D,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_1_CM8I);
  x_grlfpc2_0_comb_un1_fpci_4_2: CM8 port map (
      D0 => GRLFPC2_0_COMB_UN1_FPCI_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2_CM8I,
      S01 => GRLFPC2_0_R_A_RS2(0),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_2);
  x_grlfpc2_0_comb_un1_fpci_4_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_A_RS2D,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_2_CM8I);
  x_grlfpc2_0_comb_un1_fpci_4_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_A_RS2D,
      Y => GRLFPC2_0_COMB_UN1_FPCI_4_CM8I);
  x_grlfpc2_0_comb_un1_mexc: CM8 port map (
      D0 => GRLFPC2_0_COMB_UN1_MEXC_1,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_I_EXC(3),
      S01 => GRLFPC2_0_R_FSR_TEM(3),
      S10 => GRLFPC2_0_COMB_MEXC_1(1),
      S11 => GRLFPC2_0_COMB_MEXC_1(2),
      Y => GRLFPC2_0_COMB_UN1_MEXC);
  x_grlfpc2_0_comb_un1_mexc_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_COMB_UN1_MEXC_1_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_I_EXC(0),
      S01 => GRLFPC2_0_R_FSR_TEM(0),
      S10 => GRLFPC2_0_R_FSR_TEM(4),
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_MEXC_1);
  x_grlfpc2_0_comb_un1_mexc_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_I_EXC(4),
      Y => GRLFPC2_0_COMB_UN1_MEXC_1_CM8I);
  x_grlfpc2_0_comb_un1_r_a_rs1_1: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS1(0),
      D3 => GRLFPC2_0_R_A_ST,
      S00 => GRLFPC2_0_R_A_RS1D,
      S01 => NN_4,
      S10 => cpi_a_cnt(1),
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_R_A_RS1_1);
  x_grlfpc2_0_comb_un1_r_a_rs1_1_0: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS1(0),
      D3 => GRLFPC2_0_R_A_ST,
      S00 => GRLFPC2_0_R_A_RS1D,
      S01 => NN_4,
      S10 => cpi_a_cnt(1),
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0);
  x_grlfpc2_0_comb_un1_r_a_rs1_1_1: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS1(0),
      D3 => GRLFPC2_0_R_A_ST,
      S00 => GRLFPC2_0_R_A_RS1D,
      S01 => NN_4,
      S10 => cpi_a_cnt(1),
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1);
  x_grlfpc2_0_comb_un1_r_a_rs1_1_2: CM8 port map (
      D0 => GRLFPC2_0_R_A_RS1(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_R_A_RS1(0),
      D3 => GRLFPC2_0_R_A_ST,
      S00 => GRLFPC2_0_R_A_RS1D,
      S01 => NN_4,
      S10 => cpi_a_cnt(1),
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2);
  x_grlfpc2_0_comb_un2_holdn: AND4A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN,
      B => GRLFPC2_0_R_A_MOV,
      C => GRLFPC2_0_R_A_FPOP,
      D => HOLDN_1,
      Y => GRLFPC2_0_COMB_UN2_HOLDN);
  x_grlfpc2_0_comb_un2_holdn_0: AND4A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN_0,
      B => GRLFPC2_0_R_A_MOV,
      C => GRLFPC2_0_R_A_FPOP_0,
      D => HOLDN_0,
      Y => GRLFPC2_0_COMB_UN2_HOLDN_0);
  x_grlfpc2_0_comb_un2_holdn_1: AND4A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN_0,
      B => GRLFPC2_0_R_A_MOV,
      C => GRLFPC2_0_R_A_FPOP_0,
      D => HOLDN_0,
      Y => GRLFPC2_0_COMB_UN2_HOLDN_1);
  x_grlfpc2_0_comb_un2_holdn_2: AND4A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN_0,
      B => GRLFPC2_0_R_A_MOV,
      C => GRLFPC2_0_R_A_FPOP_0,
      D => HOLDN_0,
      Y => GRLFPC2_0_COMB_UN2_HOLDN_2);
  x_grlfpc2_0_comb_un2_holdn_3: AND4A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN_0,
      B => GRLFPC2_0_R_A_MOV,
      C => GRLFPC2_0_R_A_FPOP_0,
      D => HOLDN_0,
      Y => GRLFPC2_0_COMB_UN2_HOLDN_3);
  x_grlfpc2_0_comb_un3_holdn: OR2 port map (
      A => cpi_a_trap,
      B => cpi_a_annul,
      Y => GRLFPC2_0_COMB_UN3_HOLDN);
  x_grlfpc2_0_comb_un3_holdn_0: OR2 port map (
      A => cpi_a_trap,
      B => cpi_a_annul,
      Y => GRLFPC2_0_COMB_UN3_HOLDN_0);
  x_grlfpc2_0_comb_un4_lock: CM8 port map (
      D0 => NN_4,
      D1 => CPO_EXC_INT_1,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_UN4_LOCK_CM8I,
      S01 => GRLFPC2_0_N_331,
      S10 => cpi_d_trap,
      S11 => cpi_d_annul,
      Y => GRLFPC2_0_COMB_UN4_LOCK);
  x_grlfpc2_0_comb_un4_lock_cm8i: CM8INV port map (
      A => cpi_flush,
      Y => GRLFPC2_0_COMB_UN4_LOCK_CM8I);
  x_grlfpc2_0_comb_un6_iuexec: OR3B port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0,
      B => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK,
      C => GRLFPC2_0_COMB_UN10_IUEXEC,
      Y => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_comb_un6_iuexec_0: AND2A port map (
      A => GRLFPC2_0_R_MK_BUSY,
      B => GRLFPC2_0_R_MK_BUSY2,
      Y => GRLFPC2_0_COMB_UN6_IUEXEC_0);
  x_grlfpc2_0_comb_un6_iuexec_0_0: OR3B port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0,
      B => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK,
      C => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      Y => GRLFPC2_0_COMB_UN6_IUEXEC_0_0);
  x_grlfpc2_0_comb_un6_iuexec_1: OR3B port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0,
      B => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK,
      C => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      Y => GRLFPC2_0_COMB_UN6_IUEXEC_1);
  x_grlfpc2_0_comb_un6_iuexec_2: OR3B port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0,
      B => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK,
      C => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      Y => GRLFPC2_0_COMB_UN6_IUEXEC_2);
  x_grlfpc2_0_comb_un6_iuexec_3: OR3B port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0,
      B => GRLFPC2_0_COMB_LOCKGEN_DEPCHECK,
      C => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      Y => GRLFPC2_0_COMB_UN6_IUEXEC_3);
  x_grlfpc2_0_comb_un8_ccv: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => cpi_x_inst(19),
      S01 => GRLFPC2_0_R_X_FPOP,
      S10 => GRLFPC2_0_COMB_UN8_CCV_1,
      S11 => GRLFPC2_0_COMB_UN9_CCV,
      Y => cpo_ccv);
  x_grlfpc2_0_comb_un8_ccv_1: CM8 port map (
      D0 => GRLFPC2_0_R_E_FPOP,
      D1 => NN_4,
      D2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA,
      D3 => NN_4,
      S00 => cpi_m_inst(19),
      S01 => GRLFPC2_0_R_M_FPOP,
      S10 => GRLFPC2_0_COMB_UN8_CCV_1_CM8I,
      S11 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA,
      Y => GRLFPC2_0_COMB_UN8_CCV_1);
  x_grlfpc2_0_comb_un8_ccv_1_cm8i: CM8INV port map (
      A => cpi_e_inst(19),
      Y => GRLFPC2_0_COMB_UN8_CCV_1_CM8I);
  x_grlfpc2_0_comb_un9_ccv: AND2 port map (
      A => GRLFPC2_0_R_I_EXEC,
      B => GRLFPC2_0_R_I_INST(19),
      Y => GRLFPC2_0_COMB_UN9_CCV);
  x_grlfpc2_0_comb_un10_iuexec: OR2 port map (
      A => GRLFPC2_0_R_MK_RST2,
      B => GRLFPC2_0_R_MK_RST,
      Y => GRLFPC2_0_COMB_UN10_IUEXEC);
  x_grlfpc2_0_comb_un10_iuexec_0: OR2 port map (
      A => GRLFPC2_0_R_MK_RST2,
      B => GRLFPC2_0_R_MK_RST,
      Y => GRLFPC2_0_COMB_UN10_IUEXEC_0);
  x_grlfpc2_0_comb_v_a_afq_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_AFQ3_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_A_AFQ_1_CM8I,
      S01 => GRLFPC2_0_COMB_V_A_AFQ_1_1_0,
      S10 => cpi_d_inst(23),
      S11 => GRLFPC2_0_COMB_UN4_LOCK,
      Y => GRLFPC2_0_COMB_V_A_AFQ_1);
  x_grlfpc2_0_comb_v_a_afq_1_1_0: AND2 port map (
      A => GRLFPC2_0_COMB_RDD_1_1,
      B => GRLFPC2_0_COMB_FPDECODE_AFQ13,
      Y => GRLFPC2_0_COMB_V_A_AFQ_1_1_0);
  x_grlfpc2_0_comb_v_a_afq_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_N_17_1,
      Y => GRLFPC2_0_COMB_V_A_AFQ_1_CM8I);
  x_grlfpc2_0_comb_v_a_afsr_1: AND4B port map (
      A => GRLFPC2_0_COMB_UN4_LOCK,
      B => cpi_d_inst(20),
      C => GRLFPC2_0_N_17_1,
      D => GRLFPC2_0_COMB_V_A_AFQ_1_1_0,
      Y => GRLFPC2_0_COMB_V_A_AFSR_1);
  x_grlfpc2_0_comb_v_a_ld_1: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_A_LD_1_CM8I,
      S01 => GRLFPC2_0_COMB_FPDECODE_AFQ6_N,
      S10 => GRLFPC2_0_COMB_UN4_LOCK,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_A_LD_1);
  x_grlfpc2_0_comb_v_a_ld_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_SEQERR_UN11_OP_0,
      Y => GRLFPC2_0_COMB_V_A_LD_1_CM8I);
  x_grlfpc2_0_comb_v_a_seqerr_1: CM8 port map (
      D0 => GRLFPC2_0_COMB_V_A_AFQ_1,
      D1 => NN_2,
      D2 => GRLFPC2_0_COMB_SEQERR_UN7_OP,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN4_LOCK,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_QNE2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_A_SEQERR_1);
  x_grlfpc2_0_comb_v_a_st_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN4_LOCK,
      B => GRLFPC2_0_COMB_FPDECODE_ST,
      Y => GRLFPC2_0_COMB_V_A_ST_1);
  x_grlfpc2_0_comb_v_e_afq_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN,
      B => GRLFPC2_0_R_A_AFQ_0,
      Y => GRLFPC2_0_COMB_V_E_AFQ_1);
  x_grlfpc2_0_comb_v_e_afsr_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN,
      B => GRLFPC2_0_R_A_AFSR_0,
      Y => GRLFPC2_0_COMB_V_E_AFSR_1);
  x_grlfpc2_0_comb_v_e_fpop_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN,
      B => GRLFPC2_0_R_A_FPOP,
      Y => GRLFPC2_0_COMB_V_E_FPOP_1);
  x_grlfpc2_0_comb_v_e_ld_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN3_HOLDN,
      B => GRLFPC2_0_R_A_LD,
      Y => GRLFPC2_0_COMB_V_E_LD_1);
  x_grlfpc2_0_comb_v_e_stdata2: AND2A port map (
      A => cpi_a_cnt(1),
      B => cpi_a_cnt(0),
      Y => GRLFPC2_0_COMB_V_E_STDATA2);
  x_grlfpc2_0_comb_v_e_stdata2_0: AND2A port map (
      A => cpi_a_cnt(1),
      B => cpi_a_cnt(0),
      Y => GRLFPC2_0_COMB_V_E_STDATA2_0);
  x_grlfpc2_0_comb_v_e_stdata2_1: AND2A port map (
      A => cpi_a_cnt(1),
      B => cpi_a_cnt(0),
      Y => GRLFPC2_0_COMB_V_E_STDATA2_1);
  x_grlfpc2_0_comb_v_e_stdata2_2: AND2A port map (
      A => cpi_a_cnt(1),
      B => cpi_a_cnt(0),
      Y => GRLFPC2_0_COMB_V_E_STDATA2_2);
  x_grlfpc2_0_comb_v_e_stdata_1_0_5x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(5),
      D1 => GRLFPC2_0_R_I_PC(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_895);
  x_grlfpc2_0_comb_v_e_stdata_1_0_7x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(7),
      D1 => GRLFPC2_0_R_I_PC(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_897);
  x_grlfpc2_0_comb_v_e_stdata_1_0_8x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(8),
      D1 => GRLFPC2_0_R_I_PC(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_898);
  x_grlfpc2_0_comb_v_e_stdata_1_0_10x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(10),
      D1 => GRLFPC2_0_R_I_PC(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_900);
  x_grlfpc2_0_comb_v_e_stdata_1_0_11x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(11),
      D1 => GRLFPC2_0_R_I_PC(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_901);
  x_grlfpc2_0_comb_v_e_stdata_1_0_12x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(12),
      D1 => GRLFPC2_0_R_I_PC(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_902);
  x_grlfpc2_0_comb_v_e_stdata_1_0_13x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(13),
      D1 => GRLFPC2_0_R_I_PC(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_903);
  x_grlfpc2_0_comb_v_e_stdata_1_0_14x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(14),
      D1 => GRLFPC2_0_R_I_PC(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_904);
  x_grlfpc2_0_comb_v_e_stdata_1_0_15x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(15),
      D1 => GRLFPC2_0_R_I_PC(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_905);
  x_grlfpc2_0_comb_v_e_stdata_1_0_16x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(16),
      D1 => GRLFPC2_0_R_I_PC(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_906);
  x_grlfpc2_0_comb_v_e_stdata_1_0_17x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(17),
      D1 => GRLFPC2_0_R_I_PC(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_907);
  x_grlfpc2_0_comb_v_e_stdata_1_0_18x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(18),
      D1 => GRLFPC2_0_R_I_PC(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_908);
  x_grlfpc2_0_comb_v_e_stdata_1_0_19x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(19),
      D1 => GRLFPC2_0_R_I_PC(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_909);
  x_grlfpc2_0_comb_v_e_stdata_1_0_20x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(20),
      D1 => GRLFPC2_0_R_I_PC(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_910);
  x_grlfpc2_0_comb_v_e_stdata_1_0_21x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(21),
      D1 => GRLFPC2_0_R_I_PC(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_911);
  x_grlfpc2_0_comb_v_e_stdata_1_0_22x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(22),
      D1 => GRLFPC2_0_R_I_PC(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_912);
  x_grlfpc2_0_comb_v_e_stdata_1_0_23x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(23),
      D1 => GRLFPC2_0_R_I_PC(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_913);
  x_grlfpc2_0_comb_v_e_stdata_1_0_24x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(24),
      D1 => GRLFPC2_0_R_I_PC(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_914);
  x_grlfpc2_0_comb_v_e_stdata_1_0_25x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(25),
      D1 => GRLFPC2_0_R_I_PC(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_915);
  x_grlfpc2_0_comb_v_e_stdata_1_0_26x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(26),
      D1 => GRLFPC2_0_R_I_PC(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_916);
  x_grlfpc2_0_comb_v_e_stdata_1_0_27x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(27),
      D1 => GRLFPC2_0_R_I_PC(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_917);
  x_grlfpc2_0_comb_v_e_stdata_1_0_28x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(28),
      D1 => GRLFPC2_0_R_I_PC(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_918);
  x_grlfpc2_0_comb_v_e_stdata_1_0_29x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(29),
      D1 => GRLFPC2_0_R_I_PC(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_919);
  x_grlfpc2_0_comb_v_e_stdata_1_0_30x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(30),
      D1 => GRLFPC2_0_R_I_PC(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_920);
  x_grlfpc2_0_comb_v_e_stdata_1_1_0x: CM8 port map (
      D0 => GRLFPC2_0_OP1(32),
      D1 => GRLFPC2_0_R_FSR_CEXC(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_923);
  x_grlfpc2_0_comb_v_e_stdata_1_1_1x: CM8 port map (
      D0 => GRLFPC2_0_OP1(33),
      D1 => GRLFPC2_0_R_FSR_CEXC(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_924);
  x_grlfpc2_0_comb_v_e_stdata_1_1_2x: CM8 port map (
      D0 => GRLFPC2_0_OP1(34),
      D1 => GRLFPC2_0_R_FSR_CEXC(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_925);
  x_grlfpc2_0_comb_v_e_stdata_1_1_3x: CM8 port map (
      D0 => GRLFPC2_0_OP1(35),
      D1 => GRLFPC2_0_R_FSR_CEXC(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_926);
  x_grlfpc2_0_comb_v_e_stdata_1_1_4x: CM8 port map (
      D0 => GRLFPC2_0_OP1(36),
      D1 => GRLFPC2_0_R_FSR_CEXC(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_927);
  x_grlfpc2_0_comb_v_e_stdata_1_1_6x: CM8 port map (
      D0 => GRLFPC2_0_OP1(38),
      D1 => GRLFPC2_0_R_FSR_AEXC(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_929);
  x_grlfpc2_0_comb_v_e_stdata_1_1_9x: CM8 port map (
      D0 => GRLFPC2_0_OP1(41),
      D1 => GRLFPC2_0_R_FSR_AEXC(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_932);
  x_grlfpc2_0_comb_v_e_stdata_1_1_31x: CM8 port map (
      D0 => GRLFPC2_0_OP1(63),
      D1 => GRLFPC2_0_R_FSR_RD(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFSR_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_954);
  x_grlfpc2_0_comb_v_e_stdata_1_u_0x: CM8 port map (
      D0 => GRLFPC2_0_N_923,
      D1 => GRLFPC2_0_R_I_INST(0),
      D2 => GRLFPC2_0_N_923,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(0));
  x_grlfpc2_0_comb_v_e_stdata_1_u_1x: CM8 port map (
      D0 => GRLFPC2_0_N_924,
      D1 => GRLFPC2_0_R_I_INST(1),
      D2 => GRLFPC2_0_N_924,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(1));
  x_grlfpc2_0_comb_v_e_stdata_1_u_2x: CM8 port map (
      D0 => GRLFPC2_0_N_925,
      D1 => GRLFPC2_0_R_I_INST(2),
      D2 => GRLFPC2_0_N_925,
      D3 => GRLFPC2_0_R_I_PC(2),
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(2));
  x_grlfpc2_0_comb_v_e_stdata_1_u_3x: CM8 port map (
      D0 => GRLFPC2_0_N_926,
      D1 => GRLFPC2_0_R_I_INST(3),
      D2 => GRLFPC2_0_N_926,
      D3 => GRLFPC2_0_R_I_PC(3),
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(3));
  x_grlfpc2_0_comb_v_e_stdata_1_u_4x: CM8 port map (
      D0 => GRLFPC2_0_N_927,
      D1 => GRLFPC2_0_R_I_INST(4),
      D2 => GRLFPC2_0_N_927,
      D3 => GRLFPC2_0_R_I_PC(4),
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(4));
  x_grlfpc2_0_comb_v_e_stdata_1_u_5x: CM8 port map (
      D0 => GRLFPC2_0_OP1(37),
      D1 => GRLFPC2_0_N_895,
      D2 => GRLFPC2_0_R_FSR_AEXC(0),
      D3 => GRLFPC2_0_N_895,
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(5));
  x_grlfpc2_0_comb_v_e_stdata_1_u_6x: CM8 port map (
      D0 => GRLFPC2_0_N_929,
      D1 => GRLFPC2_0_R_I_INST(6),
      D2 => GRLFPC2_0_N_929,
      D3 => GRLFPC2_0_R_I_PC(6),
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(6));
  x_grlfpc2_0_comb_v_e_stdata_1_u_7x: CM8 port map (
      D0 => GRLFPC2_0_OP1(39),
      D1 => GRLFPC2_0_N_897,
      D2 => GRLFPC2_0_R_FSR_AEXC(2),
      D3 => GRLFPC2_0_N_897,
      S00 => GRLFPC2_0_R_A_AFQ_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(7));
  x_grlfpc2_0_comb_v_e_stdata_1_u_8x: CM8 port map (
      D0 => GRLFPC2_0_OP1(40),
      D1 => GRLFPC2_0_N_898,
      D2 => GRLFPC2_0_R_FSR_AEXC(3),
      D3 => GRLFPC2_0_N_898,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(8));
  x_grlfpc2_0_comb_v_e_stdata_1_u_9x: CM8 port map (
      D0 => GRLFPC2_0_N_932,
      D1 => GRLFPC2_0_R_I_INST(9),
      D2 => GRLFPC2_0_N_932,
      D3 => GRLFPC2_0_R_I_PC(9),
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(9));
  x_grlfpc2_0_comb_v_e_stdata_1_u_10x: CM8 port map (
      D0 => GRLFPC2_0_OP1(42),
      D1 => GRLFPC2_0_N_900,
      D2 => CPO_CC_0_INT_2,
      D3 => GRLFPC2_0_N_900,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(10));
  x_grlfpc2_0_comb_v_e_stdata_1_u_11x: CM8 port map (
      D0 => GRLFPC2_0_OP1(43),
      D1 => GRLFPC2_0_N_901,
      D2 => CPO_CC_1_INT_3,
      D3 => GRLFPC2_0_N_901,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(11));
  x_grlfpc2_0_comb_v_e_stdata_1_u_12x: CM8 port map (
      D0 => GRLFPC2_0_OP1(44),
      D1 => GRLFPC2_0_N_902,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_902,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(12));
  x_grlfpc2_0_comb_v_e_stdata_1_u_13x: CM8 port map (
      D0 => GRLFPC2_0_OP1(45),
      D1 => GRLFPC2_0_N_903,
      D2 => GRLFPC2_0_COMB_QNE2,
      D3 => GRLFPC2_0_N_903,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(13));
  x_grlfpc2_0_comb_v_e_stdata_1_u_14x: CM8 port map (
      D0 => GRLFPC2_0_OP1(46),
      D1 => GRLFPC2_0_N_904,
      D2 => GRLFPC2_0_R_FSR_FTT(0),
      D3 => GRLFPC2_0_N_904,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(14));
  x_grlfpc2_0_comb_v_e_stdata_1_u_15x: CM8 port map (
      D0 => GRLFPC2_0_OP1(47),
      D1 => GRLFPC2_0_N_905,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_905,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(15));
  x_grlfpc2_0_comb_v_e_stdata_1_u_16x: CM8 port map (
      D0 => GRLFPC2_0_OP1(48),
      D1 => GRLFPC2_0_N_906,
      D2 => GRLFPC2_0_R_FSR_FTT(2),
      D3 => GRLFPC2_0_N_906,
      S00 => GRLFPC2_0_R_A_AFQ_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(16));
  x_grlfpc2_0_comb_v_e_stdata_1_u_17x: CM8 port map (
      D0 => GRLFPC2_0_OP1(49),
      D1 => GRLFPC2_0_N_907,
      D2 => NN_4,
      D3 => GRLFPC2_0_N_907,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(17));
  x_grlfpc2_0_comb_v_e_stdata_1_u_18x: CM8 port map (
      D0 => GRLFPC2_0_OP1(50),
      D1 => GRLFPC2_0_N_908,
      D2 => NN_4,
      D3 => GRLFPC2_0_N_908,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(18));
  x_grlfpc2_0_comb_v_e_stdata_1_u_19x: CM8 port map (
      D0 => GRLFPC2_0_OP1(51),
      D1 => GRLFPC2_0_N_909,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_909,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(19));
  x_grlfpc2_0_comb_v_e_stdata_1_u_20x: CM8 port map (
      D0 => GRLFPC2_0_OP1(52),
      D1 => GRLFPC2_0_N_910,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_910,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(20));
  x_grlfpc2_0_comb_v_e_stdata_1_u_21x: CM8 port map (
      D0 => GRLFPC2_0_OP1(53),
      D1 => GRLFPC2_0_N_911,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_911,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(21));
  x_grlfpc2_0_comb_v_e_stdata_1_u_22x: CM8 port map (
      D0 => GRLFPC2_0_OP1(54),
      D1 => GRLFPC2_0_N_912,
      D2 => GRLFPC2_0_R_FSR_NONSTD,
      D3 => GRLFPC2_0_N_912,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(22));
  x_grlfpc2_0_comb_v_e_stdata_1_u_23x: CM8 port map (
      D0 => GRLFPC2_0_OP1(55),
      D1 => GRLFPC2_0_N_913,
      D2 => GRLFPC2_0_R_FSR_TEM(0),
      D3 => GRLFPC2_0_N_913,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(23));
  x_grlfpc2_0_comb_v_e_stdata_1_u_24x: CM8 port map (
      D0 => GRLFPC2_0_OP1(56),
      D1 => GRLFPC2_0_N_914,
      D2 => GRLFPC2_0_R_FSR_TEM(1),
      D3 => GRLFPC2_0_N_914,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(24));
  x_grlfpc2_0_comb_v_e_stdata_1_u_25x: CM8 port map (
      D0 => GRLFPC2_0_OP1(57),
      D1 => GRLFPC2_0_N_915,
      D2 => GRLFPC2_0_R_FSR_TEM(2),
      D3 => GRLFPC2_0_N_915,
      S00 => GRLFPC2_0_R_A_AFQ_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(25));
  x_grlfpc2_0_comb_v_e_stdata_1_u_26x: CM8 port map (
      D0 => GRLFPC2_0_OP1(58),
      D1 => GRLFPC2_0_N_916,
      D2 => GRLFPC2_0_R_FSR_TEM(3),
      D3 => GRLFPC2_0_N_916,
      S00 => GRLFPC2_0_R_A_AFQ,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(26));
  x_grlfpc2_0_comb_v_e_stdata_1_u_27x: CM8 port map (
      D0 => GRLFPC2_0_OP1(59),
      D1 => GRLFPC2_0_N_917,
      D2 => GRLFPC2_0_R_FSR_TEM(4),
      D3 => GRLFPC2_0_N_917,
      S00 => GRLFPC2_0_R_A_AFQ,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(27));
  x_grlfpc2_0_comb_v_e_stdata_1_u_28x: CM8 port map (
      D0 => GRLFPC2_0_OP1(60),
      D1 => GRLFPC2_0_N_918,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_918,
      S00 => GRLFPC2_0_R_A_AFQ,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(28));
  x_grlfpc2_0_comb_v_e_stdata_1_u_29x: CM8 port map (
      D0 => GRLFPC2_0_OP1(61),
      D1 => GRLFPC2_0_N_919,
      D2 => NN_2,
      D3 => GRLFPC2_0_N_919,
      S00 => GRLFPC2_0_R_A_AFQ,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(29));
  x_grlfpc2_0_comb_v_e_stdata_1_u_30x: CM8 port map (
      D0 => GRLFPC2_0_OP1(62),
      D1 => GRLFPC2_0_N_920,
      D2 => GRLFPC2_0_R_FSR_RD(0),
      D3 => GRLFPC2_0_N_920,
      S00 => GRLFPC2_0_R_A_AFQ,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_A_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(30));
  x_grlfpc2_0_comb_v_e_stdata_1_u_31x: CM8 port map (
      D0 => GRLFPC2_0_N_954,
      D1 => GRLFPC2_0_R_I_INST(31),
      D2 => GRLFPC2_0_N_954,
      D3 => GRLFPC2_0_R_I_PC(31),
      S00 => GRLFPC2_0_R_A_AFQ,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_V_E_STDATA2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_E_STDATA_1(31));
  x_grlfpc2_0_comb_v_fsr_aexc_1_0_0x: CM8 port map (
      D0 => GRLFPC2_0_R_FSR_AEXC(0),
      D1 => NN_4,
      D2 => cpi_dbg_data(5),
      D3 => cpi_dbg_data(5),
      S00 => GRLFPC2_0_R_I_EXC(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_664);
  x_grlfpc2_0_comb_v_fsr_aexc_1_0_1x: CM8 port map (
      D0 => GRLFPC2_0_R_FSR_AEXC(1),
      D1 => NN_4,
      D2 => cpi_dbg_data(6),
      D3 => cpi_dbg_data(6),
      S00 => GRLFPC2_0_R_I_EXC(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_665);
  x_grlfpc2_0_comb_v_fsr_aexc_1_0_2x: CM8 port map (
      D0 => GRLFPC2_0_R_FSR_AEXC(2),
      D1 => NN_4,
      D2 => cpi_dbg_data(7),
      D3 => cpi_dbg_data(7),
      S00 => GRLFPC2_0_R_I_EXC(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_666);
  x_grlfpc2_0_comb_v_fsr_aexc_1_0_3x: CM8 port map (
      D0 => GRLFPC2_0_R_FSR_AEXC(3),
      D1 => NN_4,
      D2 => cpi_dbg_data(8),
      D3 => cpi_dbg_data(8),
      S00 => GRLFPC2_0_R_I_EXC(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_667);
  x_grlfpc2_0_comb_v_fsr_aexc_1_0_4x: CM8 port map (
      D0 => GRLFPC2_0_R_FSR_AEXC(4),
      D1 => NN_4,
      D2 => cpi_dbg_data(9),
      D3 => cpi_dbg_data(9),
      S00 => GRLFPC2_0_R_I_EXC(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_668);
  x_grlfpc2_0_comb_v_fsr_aexc_1_sn_m3: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1,
      S01 => GRLFPC2_0_COMB_CCWR4_1,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => GRLFPC2_0_COMB_WRRES4,
      Y => GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4);
  x_grlfpc2_0_comb_v_fsr_aexc_1_sn_m3_436: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1,
      S01 => GRLFPC2_0_COMB_CCWR4_1,
      S10 => GRLFPC2_0_COMB_WRRES4,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1063_3);
  x_grlfpc2_0_comb_v_fsr_aexc_1_u_0x: CM8 port map (
      D0 => GRLFPC2_0_N_664,
      D1 => GRLFPC2_0_R_FSR_AEXC(0),
      D2 => GRLFPC2_0_N_664,
      D3 => cpi_lddata(5),
      S00 => GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_AEXC_1(0));
  x_grlfpc2_0_comb_v_fsr_aexc_1_u_1x: CM8 port map (
      D0 => GRLFPC2_0_N_665,
      D1 => GRLFPC2_0_R_FSR_AEXC(1),
      D2 => GRLFPC2_0_N_665,
      D3 => cpi_lddata(6),
      S00 => GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_AEXC_1(1));
  x_grlfpc2_0_comb_v_fsr_aexc_1_u_2x: CM8 port map (
      D0 => GRLFPC2_0_N_666,
      D1 => GRLFPC2_0_R_FSR_AEXC(2),
      D2 => GRLFPC2_0_N_666,
      D3 => cpi_lddata(7),
      S00 => GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_AEXC_1(2));
  x_grlfpc2_0_comb_v_fsr_aexc_1_u_3x: CM8 port map (
      D0 => GRLFPC2_0_N_667,
      D1 => GRLFPC2_0_R_FSR_AEXC(3),
      D2 => GRLFPC2_0_N_667,
      D3 => cpi_lddata(8),
      S00 => GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_AEXC_1(3));
  x_grlfpc2_0_comb_v_fsr_aexc_1_u_4x: CM8 port map (
      D0 => GRLFPC2_0_N_668,
      D1 => GRLFPC2_0_R_FSR_AEXC(4),
      D2 => GRLFPC2_0_N_668,
      D3 => cpi_lddata(9),
      S00 => GRLFPC2_0_COMB_V_FSR_AEXC_1_SN_N_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_AEXC_1(4));
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_0x: CM8 port map (
      D0 => NN_2,
      D1 => cpi_dbg_data(0),
      D2 => GRLFPC2_0_R_I_EXC(0),
      D3 => cpi_dbg_data(0),
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S01 => GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I(0),
      S10 => GRLFPC2_0_R_FSR_TEM(0),
      S11 => GRLFPC2_0_N_640,
      Y => GRLFPC2_0_N_642);
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_1x: CM8 port map (
      D0 => GRLFPC2_0_COMB_MEXC_1(1),
      D1 => GRLFPC2_0_R_I_EXC(1),
      D2 => cpi_dbg_data(1),
      D3 => GRLFPC2_0_R_I_EXC(1),
      S00 => GRLFPC2_0_N_640,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_643);
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_2x: CM8 port map (
      D0 => GRLFPC2_0_COMB_MEXC_1(2),
      D1 => GRLFPC2_0_R_I_EXC(2),
      D2 => cpi_dbg_data(2),
      D3 => GRLFPC2_0_R_I_EXC(2),
      S00 => GRLFPC2_0_N_640,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_644);
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_3x: CM8 port map (
      D0 => NN_2,
      D1 => cpi_dbg_data(3),
      D2 => GRLFPC2_0_R_I_EXC(3),
      D3 => cpi_dbg_data(3),
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      S01 => GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I(3),
      S10 => GRLFPC2_0_R_FSR_TEM(3),
      S11 => GRLFPC2_0_N_640,
      Y => GRLFPC2_0_N_645);
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_4x: CM8 port map (
      D0 => NN_2,
      D1 => cpi_dbg_data(4),
      D2 => GRLFPC2_0_R_I_EXC(4),
      D3 => cpi_dbg_data(4),
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      S01 => GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I(4),
      S10 => GRLFPC2_0_R_FSR_TEM(4),
      S11 => GRLFPC2_0_N_640,
      Y => GRLFPC2_0_N_646);
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_N_640,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I(0));
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_N_640,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I(3));
  x_grlfpc2_0_comb_v_fsr_cexc_1_2_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_N_640,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1_2_CM8I(4));
  x_grlfpc2_0_comb_v_fsr_cexc_1_sn_m2: AND2B port map (
      A => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      B => GRLFPC2_0_COMB_V_I_V6,
      Y => GRLFPC2_0_N_640);
  x_grlfpc2_0_comb_v_fsr_cexc_1_sn_m4: CM8 port map (
      D0 => GRLFPC2_0_N_640,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1,
      S01 => GRLFPC2_0_COMB_CCWR4_1,
      S10 => GRLFPC2_0_COMB_WRRES4,
      S11 => NN_2,
      Y => GRLFPC2_0_N_647);
  x_grlfpc2_0_comb_v_fsr_cexc_1_u_0x: CM8 port map (
      D0 => GRLFPC2_0_N_642,
      D1 => GRLFPC2_0_R_FSR_CEXC(0),
      D2 => GRLFPC2_0_N_642,
      D3 => cpi_lddata(0),
      S00 => GRLFPC2_0_N_647,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1(0));
  x_grlfpc2_0_comb_v_fsr_cexc_1_u_1x: CM8 port map (
      D0 => GRLFPC2_0_N_643,
      D1 => GRLFPC2_0_R_FSR_CEXC(1),
      D2 => GRLFPC2_0_N_643,
      D3 => cpi_lddata(1),
      S00 => GRLFPC2_0_N_647,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1(1));
  x_grlfpc2_0_comb_v_fsr_cexc_1_u_2x: CM8 port map (
      D0 => GRLFPC2_0_N_644,
      D1 => GRLFPC2_0_R_FSR_CEXC(2),
      D2 => GRLFPC2_0_N_644,
      D3 => cpi_lddata(2),
      S00 => GRLFPC2_0_N_647,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1(2));
  x_grlfpc2_0_comb_v_fsr_cexc_1_u_3x: CM8 port map (
      D0 => GRLFPC2_0_N_645,
      D1 => GRLFPC2_0_R_FSR_CEXC(3),
      D2 => GRLFPC2_0_N_645,
      D3 => cpi_lddata(3),
      S00 => GRLFPC2_0_N_647,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1(3));
  x_grlfpc2_0_comb_v_fsr_cexc_1_u_4x: CM8 port map (
      D0 => GRLFPC2_0_N_646,
      D1 => GRLFPC2_0_R_FSR_CEXC(4),
      D2 => GRLFPC2_0_N_646,
      D3 => cpi_lddata(4),
      S00 => GRLFPC2_0_N_647,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_CEXC_1(4));
  x_grlfpc2_0_comb_v_fsr_fcc_1_0_0x: CM8 port map (
      D0 => GRLFPC2_0_R_I_CC(0),
      D1 => cpi_dbg_data(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_655);
  x_grlfpc2_0_comb_v_fsr_fcc_1_0_1x: CM8 port map (
      D0 => GRLFPC2_0_R_I_CC(1),
      D1 => cpi_dbg_data(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_656);
  x_grlfpc2_0_comb_v_fsr_fcc_1_1_0x: CM8 port map (
      D0 => CPO_CC_0_INT_2,
      D1 => cpi_lddata(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_658);
  x_grlfpc2_0_comb_v_fsr_fcc_1_1_1x: CM8 port map (
      D0 => CPO_CC_1_INT_3,
      D1 => cpi_lddata(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_659);
  x_grlfpc2_0_comb_v_fsr_fcc_1_u_0x: CM8 port map (
      D0 => GRLFPC2_0_N_658,
      D1 => GRLFPC2_0_N_655,
      D2 => GRLFPC2_0_N_655,
      D3 => GRLFPC2_0_N_655,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1,
      S01 => GRLFPC2_0_COMB_CCWR4_1,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_FCC_1(0));
  x_grlfpc2_0_comb_v_fsr_fcc_1_u_1x: CM8 port map (
      D0 => GRLFPC2_0_N_659,
      D1 => GRLFPC2_0_N_656,
      D2 => GRLFPC2_0_N_656,
      D3 => GRLFPC2_0_N_656,
      S00 => GRLFPC2_0_COMB_ISFPOP2_1,
      S01 => GRLFPC2_0_COMB_CCWR4_1,
      S10 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_FCC_1(1));
  x_grlfpc2_0_comb_v_fsr_nonstd_1_1: AND2 port map (
      A => rst,
      B => cpi_dbg_data(22),
      Y => GRLFPC2_0_N_857);
  x_grlfpc2_0_comb_v_fsr_nonstd_1_u: CM8 port map (
      D0 => GRLFPC2_0_N_857,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_NONSTD,
      D3 => cpi_lddata(22),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_NONSTD_1);
  x_grlfpc2_0_comb_v_fsr_rd_1_1_0x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(30),
      Y => GRLFPC2_0_N_865);
  x_grlfpc2_0_comb_v_fsr_rd_1_1_1x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(31),
      Y => GRLFPC2_0_N_866);
  x_grlfpc2_0_comb_v_fsr_rd_1_u_0x: CM8 port map (
      D0 => GRLFPC2_0_N_865,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_RD(0),
      D3 => cpi_lddata(30),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_RD_1(0));
  x_grlfpc2_0_comb_v_fsr_rd_1_u_1x: CM8 port map (
      D0 => GRLFPC2_0_N_866,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_RD(1),
      D3 => cpi_lddata(31),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_RD_1(1));
  x_grlfpc2_0_comb_v_fsr_tem_1_1_0x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(23),
      Y => GRLFPC2_0_N_878);
  x_grlfpc2_0_comb_v_fsr_tem_1_1_1x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(24),
      Y => GRLFPC2_0_N_879);
  x_grlfpc2_0_comb_v_fsr_tem_1_1_2x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(25),
      Y => GRLFPC2_0_N_880);
  x_grlfpc2_0_comb_v_fsr_tem_1_1_3x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(26),
      Y => GRLFPC2_0_N_881);
  x_grlfpc2_0_comb_v_fsr_tem_1_1_4x: AND2 port map (
      A => rst,
      B => cpi_dbg_data(27),
      Y => GRLFPC2_0_N_882);
  x_grlfpc2_0_comb_v_fsr_tem_1_sn_m2: AND2B port map (
      A => RST_I,
      B => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
      Y => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3);
  x_grlfpc2_0_comb_v_fsr_tem_1_u_0x: CM8 port map (
      D0 => GRLFPC2_0_N_878,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_TEM(0),
      D3 => cpi_lddata(23),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_TEM_1(0));
  x_grlfpc2_0_comb_v_fsr_tem_1_u_1x: CM8 port map (
      D0 => GRLFPC2_0_N_879,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_TEM(1),
      D3 => cpi_lddata(24),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_TEM_1(1));
  x_grlfpc2_0_comb_v_fsr_tem_1_u_2x: CM8 port map (
      D0 => GRLFPC2_0_N_880,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_TEM(2),
      D3 => cpi_lddata(25),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_TEM_1(2));
  x_grlfpc2_0_comb_v_fsr_tem_1_u_3x: CM8 port map (
      D0 => GRLFPC2_0_N_881,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_TEM(3),
      D3 => cpi_lddata(26),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_TEM_1(3));
  x_grlfpc2_0_comb_v_fsr_tem_1_u_4x: CM8 port map (
      D0 => GRLFPC2_0_N_882,
      D1 => NN_2,
      D2 => GRLFPC2_0_R_FSR_TEM(4),
      D3 => cpi_lddata(27),
      S00 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S01 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2,
      S10 => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_FSR_TEM_1(4));
  x_grlfpc2_0_comb_v_i_exec_4: CM8 port map (
      D0 => GRLFPC2_0_R_X_FPOP,
      D1 => NN_4,
      D2 => GRLFPC2_0_R_I_EXEC,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_V_I_EXEC_4_CM8I,
      S01 => GRLFPC2_0_R_I_EXEC,
      S10 => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_EXEC_4);
  x_grlfpc2_0_comb_v_i_exec_4_cm8i: CM8INV port map (
      A => GRLFPC2_0_R_X_SEQERR,
      Y => GRLFPC2_0_COMB_V_I_EXEC_4_CM8I);
  x_grlfpc2_0_comb_v_i_inst_1_0x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(0),
      D1 => cpi_x_inst(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(0));
  x_grlfpc2_0_comb_v_i_inst_1_1x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(1),
      D1 => cpi_x_inst(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(1));
  x_grlfpc2_0_comb_v_i_inst_1_2x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(2),
      D1 => cpi_x_inst(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(2));
  x_grlfpc2_0_comb_v_i_inst_1_3x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(3),
      D1 => cpi_x_inst(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(3));
  x_grlfpc2_0_comb_v_i_inst_1_4x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(4),
      D1 => cpi_x_inst(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(4));
  x_grlfpc2_0_comb_v_i_inst_1_5x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(5),
      D1 => cpi_x_inst(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(5));
  x_grlfpc2_0_comb_v_i_inst_1_6x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(6),
      D1 => cpi_x_inst(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(6));
  x_grlfpc2_0_comb_v_i_inst_1_7x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(7),
      D1 => cpi_x_inst(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(7));
  x_grlfpc2_0_comb_v_i_inst_1_8x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(8),
      D1 => cpi_x_inst(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(8));
  x_grlfpc2_0_comb_v_i_inst_1_9x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(9),
      D1 => cpi_x_inst(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(9));
  x_grlfpc2_0_comb_v_i_inst_1_10x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(10),
      D1 => cpi_x_inst(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(10));
  x_grlfpc2_0_comb_v_i_inst_1_11x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(11),
      D1 => cpi_x_inst(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(11));
  x_grlfpc2_0_comb_v_i_inst_1_12x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(12),
      D1 => cpi_x_inst(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(12));
  x_grlfpc2_0_comb_v_i_inst_1_13x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(13),
      D1 => cpi_x_inst(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(13));
  x_grlfpc2_0_comb_v_i_inst_1_14x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(14),
      D1 => cpi_x_inst(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(14));
  x_grlfpc2_0_comb_v_i_inst_1_15x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(15),
      D1 => cpi_x_inst(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(15));
  x_grlfpc2_0_comb_v_i_inst_1_16x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(16),
      D1 => cpi_x_inst(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(16));
  x_grlfpc2_0_comb_v_i_inst_1_17x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(17),
      D1 => cpi_x_inst(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(17));
  x_grlfpc2_0_comb_v_i_inst_1_18x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(18),
      D1 => cpi_x_inst(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(18));
  x_grlfpc2_0_comb_v_i_inst_1_19x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(19),
      D1 => cpi_x_inst(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(19));
  x_grlfpc2_0_comb_v_i_inst_1_20x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(20),
      D1 => cpi_x_inst(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(20));
  x_grlfpc2_0_comb_v_i_inst_1_21x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(21),
      D1 => cpi_x_inst(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(21));
  x_grlfpc2_0_comb_v_i_inst_1_22x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(22),
      D1 => cpi_x_inst(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(22));
  x_grlfpc2_0_comb_v_i_inst_1_23x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(23),
      D1 => cpi_x_inst(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(23));
  x_grlfpc2_0_comb_v_i_inst_1_24x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(24),
      D1 => cpi_x_inst(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(24));
  x_grlfpc2_0_comb_v_i_inst_1_25x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(25),
      D1 => cpi_x_inst(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(25));
  x_grlfpc2_0_comb_v_i_inst_1_26x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(26),
      D1 => cpi_x_inst(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(26));
  x_grlfpc2_0_comb_v_i_inst_1_27x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(27),
      D1 => cpi_x_inst(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(27));
  x_grlfpc2_0_comb_v_i_inst_1_28x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(28),
      D1 => cpi_x_inst(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(28));
  x_grlfpc2_0_comb_v_i_inst_1_29x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(29),
      D1 => cpi_x_inst(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(29));
  x_grlfpc2_0_comb_v_i_inst_1_30x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(30),
      D1 => cpi_x_inst(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(30));
  x_grlfpc2_0_comb_v_i_inst_1_31x: CM8 port map (
      D0 => GRLFPC2_0_R_I_INST(31),
      D1 => cpi_x_inst(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_INST_1(31));
  x_grlfpc2_0_comb_v_i_pc_1_2x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(2),
      D1 => cpi_x_pc(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(2));
  x_grlfpc2_0_comb_v_i_pc_1_3x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(3),
      D1 => cpi_x_pc(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(3));
  x_grlfpc2_0_comb_v_i_pc_1_4x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(4),
      D1 => cpi_x_pc(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(4));
  x_grlfpc2_0_comb_v_i_pc_1_5x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(5),
      D1 => cpi_x_pc(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(5));
  x_grlfpc2_0_comb_v_i_pc_1_6x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(6),
      D1 => cpi_x_pc(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(6));
  x_grlfpc2_0_comb_v_i_pc_1_7x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(7),
      D1 => cpi_x_pc(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(7));
  x_grlfpc2_0_comb_v_i_pc_1_8x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(8),
      D1 => cpi_x_pc(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(8));
  x_grlfpc2_0_comb_v_i_pc_1_9x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(9),
      D1 => cpi_x_pc(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(9));
  x_grlfpc2_0_comb_v_i_pc_1_10x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(10),
      D1 => cpi_x_pc(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(10));
  x_grlfpc2_0_comb_v_i_pc_1_11x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(11),
      D1 => cpi_x_pc(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(11));
  x_grlfpc2_0_comb_v_i_pc_1_12x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(12),
      D1 => cpi_x_pc(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(12));
  x_grlfpc2_0_comb_v_i_pc_1_13x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(13),
      D1 => cpi_x_pc(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(13));
  x_grlfpc2_0_comb_v_i_pc_1_14x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(14),
      D1 => cpi_x_pc(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(14));
  x_grlfpc2_0_comb_v_i_pc_1_15x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(15),
      D1 => cpi_x_pc(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(15));
  x_grlfpc2_0_comb_v_i_pc_1_16x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(16),
      D1 => cpi_x_pc(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(16));
  x_grlfpc2_0_comb_v_i_pc_1_17x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(17),
      D1 => cpi_x_pc(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(17));
  x_grlfpc2_0_comb_v_i_pc_1_18x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(18),
      D1 => cpi_x_pc(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(18));
  x_grlfpc2_0_comb_v_i_pc_1_19x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(19),
      D1 => cpi_x_pc(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(19));
  x_grlfpc2_0_comb_v_i_pc_1_20x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(20),
      D1 => cpi_x_pc(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(20));
  x_grlfpc2_0_comb_v_i_pc_1_21x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(21),
      D1 => cpi_x_pc(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(21));
  x_grlfpc2_0_comb_v_i_pc_1_22x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(22),
      D1 => cpi_x_pc(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(22));
  x_grlfpc2_0_comb_v_i_pc_1_23x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(23),
      D1 => cpi_x_pc(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(23));
  x_grlfpc2_0_comb_v_i_pc_1_24x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(24),
      D1 => cpi_x_pc(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(24));
  x_grlfpc2_0_comb_v_i_pc_1_25x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(25),
      D1 => cpi_x_pc(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(25));
  x_grlfpc2_0_comb_v_i_pc_1_26x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(26),
      D1 => cpi_x_pc(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(26));
  x_grlfpc2_0_comb_v_i_pc_1_27x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(27),
      D1 => cpi_x_pc(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(27));
  x_grlfpc2_0_comb_v_i_pc_1_28x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(28),
      D1 => cpi_x_pc(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(28));
  x_grlfpc2_0_comb_v_i_pc_1_29x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(29),
      D1 => cpi_x_pc(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(29));
  x_grlfpc2_0_comb_v_i_pc_1_30x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(30),
      D1 => cpi_x_pc(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(30));
  x_grlfpc2_0_comb_v_i_pc_1_31x: CM8 port map (
      D0 => GRLFPC2_0_R_I_PC(31),
      D1 => cpi_x_pc(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_EXEC_0_SQMUXA,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_PC_1(31));
  x_grlfpc2_0_comb_v_i_res_1_29x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(32),
      D1 => GRLFPC2_0_R_I_RES(29),
      D2 => GRLFPC2_0_OP2(32),
      D3 => GRLFPC2_0_OP2(32),
      S00 => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(29));
  x_grlfpc2_0_comb_v_i_res_1_30x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(30),
      D1 => GRLFPC2_0_FPO_FRAC(33),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(33),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(30));
  x_grlfpc2_0_comb_v_i_res_1_31x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(31),
      D1 => GRLFPC2_0_FPO_FRAC(34),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(34),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(31));
  x_grlfpc2_0_comb_v_i_res_1_32x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(32),
      D1 => GRLFPC2_0_FPO_FRAC(35),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(35),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(32));
  x_grlfpc2_0_comb_v_i_res_1_33x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(33),
      D1 => GRLFPC2_0_FPO_FRAC(36),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(36),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(33));
  x_grlfpc2_0_comb_v_i_res_1_34x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(34),
      D1 => GRLFPC2_0_FPO_FRAC(37),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(37),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_0,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(34));
  x_grlfpc2_0_comb_v_i_res_1_35x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(35),
      D1 => GRLFPC2_0_FPO_FRAC(38),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(38),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(35));
  x_grlfpc2_0_comb_v_i_res_1_36x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(36),
      D1 => GRLFPC2_0_FPO_FRAC(39),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(39),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(36));
  x_grlfpc2_0_comb_v_i_res_1_37x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(40),
      D1 => GRLFPC2_0_R_I_RES(37),
      D2 => GRLFPC2_0_OP2(40),
      D3 => GRLFPC2_0_OP2(40),
      S00 => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(37));
  x_grlfpc2_0_comb_v_i_res_1_38x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(38),
      D1 => GRLFPC2_0_FPO_FRAC(41),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(41),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(38));
  x_grlfpc2_0_comb_v_i_res_1_39x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(39),
      D1 => GRLFPC2_0_FPO_FRAC(42),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(42),
      S00 => GRLFPC2_0_UN1_HOLDN_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(39));
  x_grlfpc2_0_comb_v_i_res_1_40x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(40),
      D1 => GRLFPC2_0_FPO_FRAC(43),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(43),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(40));
  x_grlfpc2_0_comb_v_i_res_1_41x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(41),
      D1 => GRLFPC2_0_FPO_FRAC(44),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(44),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(41));
  x_grlfpc2_0_comb_v_i_res_1_42x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(42),
      D1 => GRLFPC2_0_FPO_FRAC(45),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(45),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(42));
  x_grlfpc2_0_comb_v_i_res_1_43x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(43),
      D1 => GRLFPC2_0_FPO_FRAC(46),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(46),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(43));
  x_grlfpc2_0_comb_v_i_res_1_44x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(44),
      D1 => GRLFPC2_0_FPO_FRAC(47),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(47),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(44));
  x_grlfpc2_0_comb_v_i_res_1_45x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(45),
      D1 => GRLFPC2_0_FPO_FRAC(48),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(48),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(45));
  x_grlfpc2_0_comb_v_i_res_1_46x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(46),
      D1 => GRLFPC2_0_FPO_FRAC(49),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(49),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(46));
  x_grlfpc2_0_comb_v_i_res_1_47x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(47),
      D1 => GRLFPC2_0_FPO_FRAC(50),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(50),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(47));
  x_grlfpc2_0_comb_v_i_res_1_48x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(48),
      D1 => GRLFPC2_0_FPO_FRAC(51),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(51),
      S00 => GRLFPC2_0_UN1_HOLDN_1_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(48));
  x_grlfpc2_0_comb_v_i_res_1_49x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(49),
      D1 => GRLFPC2_0_FPO_FRAC(52),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(52),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(49));
  x_grlfpc2_0_comb_v_i_res_1_50x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(50),
      D1 => GRLFPC2_0_FPO_FRAC(53),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(53),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(50));
  x_grlfpc2_0_comb_v_i_res_1_51x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(51),
      D1 => GRLFPC2_0_FPO_FRAC_0(54),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(54),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(51));
  x_grlfpc2_0_comb_v_i_res_1_52x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(52),
      D1 => GRLFPC2_0_FPO_EXP(0),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(55),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(52));
  x_grlfpc2_0_comb_v_i_res_1_53x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(53),
      D1 => GRLFPC2_0_FPO_EXP(1),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(56),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(53));
  x_grlfpc2_0_comb_v_i_res_1_54x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(54),
      D1 => GRLFPC2_0_FPO_EXP(2),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(57),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(54));
  x_grlfpc2_0_comb_v_i_res_1_55x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(55),
      D1 => GRLFPC2_0_FPO_EXP(3),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(58),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(55));
  x_grlfpc2_0_comb_v_i_res_1_56x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(56),
      D1 => GRLFPC2_0_FPO_EXP(4),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(59),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(56));
  x_grlfpc2_0_comb_v_i_res_1_57x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(57),
      D1 => GRLFPC2_0_FPO_EXP(5),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(60),
      S00 => GRLFPC2_0_UN1_HOLDN_1_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(57));
  x_grlfpc2_0_comb_v_i_res_1_58x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(58),
      D1 => GRLFPC2_0_FPO_EXP(6),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(61),
      S00 => GRLFPC2_0_UN1_HOLDN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(58));
  x_grlfpc2_0_comb_v_i_res_1_59x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(59),
      D1 => GRLFPC2_0_FPO_EXP(7),
      D2 => NN_2,
      D3 => GRLFPC2_0_OP2(62),
      S00 => GRLFPC2_0_UN1_HOLDN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(59));
  x_grlfpc2_0_comb_v_i_res_1_63x: CM8 port map (
      D0 => GRLFPC2_0_FPO_SIGN,
      D1 => GRLFPC2_0_R_I_RES(63),
      D2 => GRLFPC2_0_COMB_V_I_RES_6(63),
      D3 => GRLFPC2_0_COMB_V_I_RES_6(63),
      S00 => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_1(63));
  x_grlfpc2_0_comb_v_i_res_6_63x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_COMB_V_I_RES_6_CM8I(63),
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_V_I_RES_6_CM8I(63),
      S01 => GRLFPC2_0_OP2(63),
      S10 => cpi_a_inst(7),
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_RES_6(63));
  x_grlfpc2_0_comb_v_i_res_6_cm8i_63x: CM8INV port map (
      A => cpi_a_inst(8),
      Y => GRLFPC2_0_COMB_V_I_RES_6_CM8I(63));
  x_grlfpc2_0_comb_v_i_v6: AND3A port map (
      A => GRLFPC2_0_COMB_UN1_MEXC,
      B => GRLFPC2_0_COMB_V_I_EXEC_4,
      C => GRLFPC2_0_R_I_V,
      Y => GRLFPC2_0_COMB_V_I_V6);
  x_grlfpc2_0_comb_v_i_v_1: CM8 port map (
      D0 => GRLFPC2_0_UN1_HOLDN_1,
      D1 => GRLFPC2_0_COMB_V_I_V_1_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_I_V_1_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_ANNULRES_1,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_I_V_1);
  x_grlfpc2_0_comb_v_i_v_1_cm8i: CM8INV port map (
      A => HOLDN_1,
      Y => GRLFPC2_0_COMB_V_I_V_1_CM8I);
  x_grlfpc2_0_comb_v_m_afq_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_2,
      B => GRLFPC2_0_R_E_AFQ,
      Y => GRLFPC2_0_COMB_V_M_AFQ_1);
  x_grlfpc2_0_comb_v_m_afsr_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_2,
      B => GRLFPC2_0_R_E_AFSR,
      Y => GRLFPC2_0_COMB_V_M_AFSR_1);
  x_grlfpc2_0_comb_v_m_fpop_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_2,
      B => GRLFPC2_0_R_E_FPOP,
      Y => GRLFPC2_0_COMB_V_M_FPOP_1);
  x_grlfpc2_0_comb_v_m_ld_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_2,
      B => GRLFPC2_0_R_E_LD,
      Y => GRLFPC2_0_COMB_V_M_LD_1);
  x_grlfpc2_0_comb_v_mk_ldop_1: AND3B port map (
      A => GRLFPC2_0_COMB_UN4_LOCK,
      B => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      C => HOLDN_1,
      Y => GRLFPC2_0_COMB_V_MK_LDOP_1);
  x_grlfpc2_0_comb_v_mk_rst_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      S10 => GRLFPC2_0_COMB_V_MK_RST_1_3,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_V_MK_RST_1);
  x_grlfpc2_0_comb_v_mk_rst_1_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_ANNULFPU_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => HOLDN_1,
      S01 => CPO_HOLDN_INT_4,
      S10 => GRLFPC2_0_R_MK_RST,
      S11 => GRLFPC2_0_R_MK_RST2,
      Y => GRLFPC2_0_COMB_V_MK_RST_1_3);
  x_grlfpc2_0_comb_v_state12: AND3A port map (
      A => GRLFPC2_0_R_STATE(1),
      B => GRLFPC2_0_R_STATE(0),
      C => cpi_exack,
      Y => GRLFPC2_0_COMB_V_STATE12);
  x_grlfpc2_0_comb_v_state_1_0x: AND3A port map (
      A => GRLFPC2_0_COMB_V_STATE12,
      B => GRLFPC2_0_COMB_V_STATE_7(0),
      C => GRLFPC2_0_V_STATE_1_SQMUXA,
      Y => GRLFPC2_0_COMB_V_STATE_1(0));
  x_grlfpc2_0_comb_v_state_1_1x: CM8 port map (
      D0 => GRLFPC2_0_V_STATE_1_SQMUXA,
      D1 => GRLFPC2_0_R_STATE(1),
      D2 => GRLFPC2_0_V_STATE_1_SQMUXA,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_STATE_1_SQMUXA,
      S01 => GRLFPC2_0_COMB_V_STATE_1_CM8I(1),
      S10 => GRLFPC2_0_UN1_FPCI_2_N,
      S11 => GRLFPC2_0_COMB_V_I_V6,
      Y => GRLFPC2_0_COMB_V_STATE_1(1));
  x_grlfpc2_0_comb_v_state_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_COMB_V_STATE12,
      Y => GRLFPC2_0_COMB_V_STATE_1_CM8I(1));
  x_grlfpc2_0_comb_v_state_7_0x: CM8 port map (
      D0 => GRLFPC2_0_R_STATE(0),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_UN1_FPCI_2_N,
      S01 => NN_4,
      S10 => GRLFPC2_0_V_FSR_FTT_0_SQMUXA_2_1,
      S11 => GRLFPC2_0_COMB_V_I_V6,
      Y => GRLFPC2_0_COMB_V_STATE_7(0));
  x_grlfpc2_0_comb_v_x_afq_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1,
      B => GRLFPC2_0_R_M_AFQ,
      Y => GRLFPC2_0_COMB_V_X_AFQ_1);
  x_grlfpc2_0_comb_v_x_afsr_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1,
      B => GRLFPC2_0_R_M_AFSR,
      Y => GRLFPC2_0_COMB_V_X_AFSR_1);
  x_grlfpc2_0_comb_v_x_fpop_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1,
      B => GRLFPC2_0_R_M_FPOP,
      Y => GRLFPC2_0_COMB_V_X_FPOP_1);
  x_grlfpc2_0_comb_v_x_ld_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1,
      B => GRLFPC2_0_R_M_LD,
      Y => GRLFPC2_0_COMB_V_X_LD_1);
  x_grlfpc2_0_comb_wrdata_4_0x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(29),
      D1 => GRLFPC2_0_R_I_RES(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(0));
  x_grlfpc2_0_comb_wrdata_4_1x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(30),
      D1 => GRLFPC2_0_R_I_RES(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(1));
  x_grlfpc2_0_comb_wrdata_4_2x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(31),
      D1 => GRLFPC2_0_R_I_RES(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(2));
  x_grlfpc2_0_comb_wrdata_4_3x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(32),
      D1 => GRLFPC2_0_R_I_RES(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(3));
  x_grlfpc2_0_comb_wrdata_4_4x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(33),
      D1 => GRLFPC2_0_R_I_RES(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(4));
  x_grlfpc2_0_comb_wrdata_4_5x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(34),
      D1 => GRLFPC2_0_R_I_RES(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(5));
  x_grlfpc2_0_comb_wrdata_4_6x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(35),
      D1 => GRLFPC2_0_R_I_RES(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(6));
  x_grlfpc2_0_comb_wrdata_4_7x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(36),
      D1 => GRLFPC2_0_R_I_RES(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(7));
  x_grlfpc2_0_comb_wrdata_4_8x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(37),
      D1 => GRLFPC2_0_R_I_RES(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(8));
  x_grlfpc2_0_comb_wrdata_4_9x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(38),
      D1 => GRLFPC2_0_R_I_RES(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(9));
  x_grlfpc2_0_comb_wrdata_4_10x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(39),
      D1 => GRLFPC2_0_R_I_RES(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(10));
  x_grlfpc2_0_comb_wrdata_4_11x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(40),
      D1 => GRLFPC2_0_R_I_RES(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(11));
  x_grlfpc2_0_comb_wrdata_4_12x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(41),
      D1 => GRLFPC2_0_R_I_RES(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(12));
  x_grlfpc2_0_comb_wrdata_4_13x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(42),
      D1 => GRLFPC2_0_R_I_RES(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(13));
  x_grlfpc2_0_comb_wrdata_4_14x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(43),
      D1 => GRLFPC2_0_R_I_RES(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(14));
  x_grlfpc2_0_comb_wrdata_4_15x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(44),
      D1 => GRLFPC2_0_R_I_RES(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(15));
  x_grlfpc2_0_comb_wrdata_4_16x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(45),
      D1 => GRLFPC2_0_R_I_RES(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(16));
  x_grlfpc2_0_comb_wrdata_4_17x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(46),
      D1 => GRLFPC2_0_R_I_RES(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(17));
  x_grlfpc2_0_comb_wrdata_4_18x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(47),
      D1 => GRLFPC2_0_R_I_RES(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(18));
  x_grlfpc2_0_comb_wrdata_4_19x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(48),
      D1 => GRLFPC2_0_R_I_RES(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(19));
  x_grlfpc2_0_comb_wrdata_4_20x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(49),
      D1 => GRLFPC2_0_R_I_RES(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(20));
  x_grlfpc2_0_comb_wrdata_4_21x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(50),
      D1 => GRLFPC2_0_R_I_RES(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(21));
  x_grlfpc2_0_comb_wrdata_4_22x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(51),
      D1 => GRLFPC2_0_R_I_RES(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(22));
  x_grlfpc2_0_comb_wrdata_4_23x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(52),
      D1 => GRLFPC2_0_R_I_RES(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(23));
  x_grlfpc2_0_comb_wrdata_4_24x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(53),
      D1 => GRLFPC2_0_R_I_RES(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(24));
  x_grlfpc2_0_comb_wrdata_4_25x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(54),
      D1 => GRLFPC2_0_R_I_RES(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(25));
  x_grlfpc2_0_comb_wrdata_4_26x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(55),
      D1 => GRLFPC2_0_R_I_RES(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(26));
  x_grlfpc2_0_comb_wrdata_4_27x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(56),
      D1 => GRLFPC2_0_R_I_RES(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(27));
  x_grlfpc2_0_comb_wrdata_4_28x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(57),
      D1 => GRLFPC2_0_R_I_RES(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(28));
  x_grlfpc2_0_comb_wrdata_4_29x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(58),
      D1 => GRLFPC2_0_R_I_RES(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(29));
  x_grlfpc2_0_comb_wrdata_4_30x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(59),
      D1 => GRLFPC2_0_R_I_RES(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(30));
  x_grlfpc2_0_comb_wrdata_4_32x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(29),
      D1 => GRLFPC2_0_R_I_RES(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(32));
  x_grlfpc2_0_comb_wrdata_4_33x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(30),
      D1 => GRLFPC2_0_R_I_RES(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(33));
  x_grlfpc2_0_comb_wrdata_4_34x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(31),
      D1 => GRLFPC2_0_R_I_RES(34),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(34));
  x_grlfpc2_0_comb_wrdata_4_35x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(32),
      D1 => GRLFPC2_0_R_I_RES(35),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(35));
  x_grlfpc2_0_comb_wrdata_4_36x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(33),
      D1 => GRLFPC2_0_R_I_RES(36),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(36));
  x_grlfpc2_0_comb_wrdata_4_37x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(34),
      D1 => GRLFPC2_0_R_I_RES(37),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(37));
  x_grlfpc2_0_comb_wrdata_4_38x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(35),
      D1 => GRLFPC2_0_R_I_RES(38),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(38));
  x_grlfpc2_0_comb_wrdata_4_39x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(36),
      D1 => GRLFPC2_0_R_I_RES(39),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(39));
  x_grlfpc2_0_comb_wrdata_4_40x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(37),
      D1 => GRLFPC2_0_R_I_RES(40),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(40));
  x_grlfpc2_0_comb_wrdata_4_41x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(38),
      D1 => GRLFPC2_0_R_I_RES(41),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(41));
  x_grlfpc2_0_comb_wrdata_4_42x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(39),
      D1 => GRLFPC2_0_R_I_RES(42),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(42));
  x_grlfpc2_0_comb_wrdata_4_43x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(40),
      D1 => GRLFPC2_0_R_I_RES(43),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(43));
  x_grlfpc2_0_comb_wrdata_4_44x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(41),
      D1 => GRLFPC2_0_R_I_RES(44),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(44));
  x_grlfpc2_0_comb_wrdata_4_45x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(42),
      D1 => GRLFPC2_0_R_I_RES(45),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(45));
  x_grlfpc2_0_comb_wrdata_4_46x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(43),
      D1 => GRLFPC2_0_R_I_RES(46),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(46));
  x_grlfpc2_0_comb_wrdata_4_47x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(44),
      D1 => GRLFPC2_0_R_I_RES(47),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(47));
  x_grlfpc2_0_comb_wrdata_4_48x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(45),
      D1 => GRLFPC2_0_R_I_RES(48),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(48));
  x_grlfpc2_0_comb_wrdata_4_49x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(46),
      D1 => GRLFPC2_0_R_I_RES(49),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(49));
  x_grlfpc2_0_comb_wrdata_4_50x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(47),
      D1 => GRLFPC2_0_R_I_RES(50),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(50));
  x_grlfpc2_0_comb_wrdata_4_51x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(48),
      D1 => GRLFPC2_0_R_I_RES(51),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(51));
  x_grlfpc2_0_comb_wrdata_4_52x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(49),
      D1 => GRLFPC2_0_R_I_RES(52),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(52));
  x_grlfpc2_0_comb_wrdata_4_53x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(50),
      D1 => GRLFPC2_0_R_I_RES(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(53));
  x_grlfpc2_0_comb_wrdata_4_54x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(51),
      D1 => GRLFPC2_0_R_I_RES(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(54));
  x_grlfpc2_0_comb_wrdata_4_55x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(52),
      D1 => GRLFPC2_0_R_I_RES(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(55));
  x_grlfpc2_0_comb_wrdata_4_56x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(53),
      D1 => GRLFPC2_0_R_I_RES(56),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(56));
  x_grlfpc2_0_comb_wrdata_4_57x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(54),
      D1 => GRLFPC2_0_R_I_RES(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3_0_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(57));
  x_grlfpc2_0_comb_wrdata_4_58x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(55),
      D1 => GRLFPC2_0_R_I_RES(58),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(58));
  x_grlfpc2_0_comb_wrdata_4_59x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(56),
      D1 => GRLFPC2_0_R_I_RES(59),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(59));
  x_grlfpc2_0_comb_wrdata_4_60x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(57),
      D1 => GRLFPC2_0_R_I_RES(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(60));
  x_grlfpc2_0_comb_wrdata_4_61x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(58),
      D1 => GRLFPC2_0_R_I_RES(61),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(61));
  x_grlfpc2_0_comb_wrdata_4_62x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(59),
      D1 => GRLFPC2_0_R_I_RES(62),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_RDD_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WRDATA_4(62));
  x_grlfpc2_0_comb_wren1_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_WREN1_1_CM8I,
      D2 => GRLFPC2_0_COMB_WREN1_9,
      D3 => GRLFPC2_0_COMB_WREN1_1_CM8I,
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => HOLDN_1,
      S11 => NN_2,
      Y => rfi1_wren);
  x_grlfpc2_0_comb_wren1_1_cm8i: CM8INV port map (
      A => cpi_dbg_addr(0),
      Y => GRLFPC2_0_COMB_WREN1_1_CM8I);
  x_grlfpc2_0_comb_wren1_9: CM8 port map (
      D0 => GRLFPC2_0_N_552,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_WREN1_0_SQMUXA_3,
      S01 => GRLFPC2_0_N_552,
      S10 => GRLFPC2_0_COMB_WREN1_9_CM8I,
      S11 => GRLFPC2_0_WREN1_M(0),
      Y => GRLFPC2_0_COMB_WREN1_9);
  x_grlfpc2_0_comb_wren1_9_cm8i: CM8INV port map (
      A => GRLFPC2_0_WREN210_M_N(340),
      Y => GRLFPC2_0_COMB_WREN1_9_CM8I);
  x_grlfpc2_0_comb_wren2_1: CM8 port map (
      D0 => NN_2,
      D1 => cpi_dbg_addr(0),
      D2 => GRLFPC2_0_COMB_WREN2_9,
      D3 => cpi_dbg_addr(0),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => HOLDN_1,
      S11 => NN_2,
      Y => rfi2_wren);
  x_grlfpc2_0_comb_wren2_9: CM8 port map (
      D0 => GRLFPC2_0_N_548,
      D1 => GRLFPC2_0_UN1_WREN1_0_SQMUXA,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_N_552,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_COMB_WREN2_9);
  x_grlfpc2_0_comb_wren2_9s_iv: CM8 port map (
      D0 => GRLFPC2_0_WREN2_2_SQMUXA_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_WREN1_M_N(0),
      S01 => GRLFPC2_0_COMB_WRRES4,
      S10 => GRLFPC2_0_COMB_WREN2_9S_IV_CM8I,
      S11 => cpi_x_inst(20),
      Y => GRLFPC2_0_N_548);
  x_grlfpc2_0_comb_wren2_9s_iv_cm8i: CM8INV port map (
      A => GRLFPC2_0_WREN210_M_N(340),
      Y => GRLFPC2_0_COMB_WREN2_9S_IV_CM8I);
  x_grlfpc2_0_comb_wren22: AND2B port map (
      A => cpi_x_cnt(0),
      B => cpi_x_cnt(1),
      Y => GRLFPC2_0_COMB_WREN22);
  x_grlfpc2_0_comb_wrres4: AND3A port map (
      A => GRLFPC2_0_COMB_V_STATE_7(0),
      B => GRLFPC2_0_COMB_CCWR4_1_0,
      C => GRLFPC2_0_COMB_WRRES4_0,
      Y => GRLFPC2_0_COMB_WRRES4);
  x_grlfpc2_0_comb_wrres4_0: AND2B port map (
      A => GRLFPC2_0_COMB_ISFPOP2_1,
      B => GRLFPC2_0_R_X_LD_0,
      Y => GRLFPC2_0_COMB_WRRES4_0);
  x_grlfpc2_0_fpco_holdn: AND2 port map (
      A => GRLFPC2_0_R_MK_HOLDN1,
      B => GRLFPC2_0_R_MK_HOLDN2,
      Y => CPO_HOLDN_INT_4);
  x_grlfpc2_0_fpi_ldop: OR3A port map (
      A => rst,
      B => GRLFPC2_0_COMB_UN10_IUEXEC,
      C => GRLFPC2_0_R_MK_LDOP,
      Y => GRLFPC2_0_FPI_LDOP);
  x_grlfpc2_0_fpi_ldop_0: OR3A port map (
      A => rst,
      B => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      C => GRLFPC2_0_R_MK_LDOP,
      Y => GRLFPC2_0_FPI_LDOP_0);
  x_grlfpc2_0_fpi_ldop_1: OR3A port map (
      A => rst,
      B => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      C => GRLFPC2_0_R_MK_LDOP,
      Y => GRLFPC2_0_FPI_LDOP_1);
  x_grlfpc2_0_fpi_ldop_2: OR3A port map (
      A => rst,
      B => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      C => GRLFPC2_0_R_MK_LDOP,
      Y => GRLFPC2_0_FPI_LDOP_2);
  x_grlfpc2_0_fpi_ldop_3: OR3A port map (
      A => rst,
      B => GRLFPC2_0_COMB_UN10_IUEXEC_0,
      C => GRLFPC2_0_R_MK_LDOP,
      Y => GRLFPC2_0_FPI_LDOP_3);
  x_grlfpc2_0_fpi_start: AND4C port map (
      A => GRLFPC2_0_COMB_UN4_LOCK,
      B => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      C => GRLFPC2_0_COMB_UN10_IUEXEC,
      D => HOLDN_1,
      Y => GRLFPC2_0_FPI_START);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_ConditionCodes_1_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONCODES_1_CM8I(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      S11 => NN_2,
      Y => GRLFPC2_0_FPO_CC(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_ConditionCodes_1_1x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONCODES_1_CM8I(1),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      S11 => NN_2,
      Y => GRLFPC2_0_FPO_CC(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_ConditionCodes_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONCODES_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_ConditionCodes_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONCODES_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_0x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_CM8I(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_26,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_27,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_0_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT,
      Y => GRLFPC2_0_FPO_EXC(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_1x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(41),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      Y => GRLFPC2_0_FPO_EXC(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_3x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      Y => GRLFPC2_0_FPO_EXC(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_4x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(41),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      S11 => NN_2,
      Y => GRLFPC2_0_FPO_EXC(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_0_2x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_25,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1766_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1766_N_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1766_N_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3275_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1766_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1766_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1768: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1768_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1768_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3277);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1768_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1768_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1769: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1769_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1769_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3713,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3278);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1769_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1769_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1770: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1770_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1770_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3714,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3279);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1770_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1770_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1773: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1773_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1773_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3717,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3282);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1773_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1773_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1777: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(12),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3286);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1783_n: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3310_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1785: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3312);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1786: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1786_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1786_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3313_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1786_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1786_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1787: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1787_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1787_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3314_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1787_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1787_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1789: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1789_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1789_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3316_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1789_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1789_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1791: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1791_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1791_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3318);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1791_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1791_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1792: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1792_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1792_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3319);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1792_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1792_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1795: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1795_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1795_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3322_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1795_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1795_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1796_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1796_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1797: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1797_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1797_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3324);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1797_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1797_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1798: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(15),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3325);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1799: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1799_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1799_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3326);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1799_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1799_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1800: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1800_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1800_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3327);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1800_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1800_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1802: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1802_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1802_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(19),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3329);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1802_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1802_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1803: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(20),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3330);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1804: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1804_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1804_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(21),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3331);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1804_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1804_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1806: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1806_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1806_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(23),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3333);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1806_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1806_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1807: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1807_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1807_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(24),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3334_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1807_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1807_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1808: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1808_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1808_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(25),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3335_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1808_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1808_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1811: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1811_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1811_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(28),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3338_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1811_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1811_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1812_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1812_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1813: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(30),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3340);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1815: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1815_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1815_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(32),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3342);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1815_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1815_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1816: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1816_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1816_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(33),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3343);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1816_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1816_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1819: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(36),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3346);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1820: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(37),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3347);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1821: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(38),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1821_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1821_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(38),
      S01 => NN_4,
      S10 => NN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3348);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1821_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1821_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1823: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(40),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1823_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1823_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3350);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1823_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1823_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1824: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1824_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1824_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3351);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1824_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1824_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1828_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1828_N_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1828_N_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3355_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1828_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1828_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1829: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(46),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3356);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1830_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1830_N_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1830_N_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3357_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1830_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1830_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1831_s: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(48),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1831_s_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1833: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(50),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3360);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1836_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1836_N_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1836_N_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3363_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1836_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1836_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1838: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1838_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1838_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(55),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3365_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_1838_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1838_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_SignResult: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SIGNRESULT_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN1_GRFPUS,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(23),
      S11 => NN_2,
      Y => GRLFPC2_0_FPO_SIGN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_SignResult_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SIGNRESULT_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un5_notainfnan: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      S10 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un5_notainfnan_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un5_notazerodenorm: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(236),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(235),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un5_notbzerodenorm_n: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un11_notbinfnan_n: OR3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTBINFNAN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notainfnan_4_n: OR4D port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notainfnan_5: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notainfnan_n: OR3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notbinfnan_0: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notbinfnan_4: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notbinfnan_6_n: OR4D port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_4,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_6_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_busymulxff_un2_temp_1: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(70),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_busymulxff_un2_temp_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_busymulxff_un2_temp_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_checkovanddenorm_un20_notpossibleov: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_FPO_FRAC_0(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_FPO_FRAC(53),
      S01 => GRLFPC2_0_FPO_FRAC(52),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_4_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_checkovanddenorm_un20_notpossibleov_4_n: OR4D port map (
      A => GRLFPC2_0_FPO_FRAC(51),
      B => GRLFPC2_0_FPO_FRAC(50),
      C => GRLFPC2_0_FPO_FRAC(48),
      D => GRLFPC2_0_FPO_FRAC(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_4_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_checkovanddenorm_un20_notpossibleov_cm8i: CM8INV port map (
      A => GRLFPC2_0_FPO_FRAC(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_condmuxmulxff_un4_notsqrtlftcc: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpAregLC_0x: AND2A port map (
      A => GRLFPC2_0_FPI_LDOP_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpAregLoadEn: CM8 port map (
      D0 => GRLFPC2_0_FPI_LDOP_0,
      D1 => GRLFPC2_0_FPI_LDOP_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_CM8I,
      D3 => GRLFPC2_0_FPI_LDOP_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpAregLoadEn_0: CM8 port map (
      D0 => GRLFPC2_0_FPI_LDOP_0,
      D1 => GRLFPC2_0_FPI_LDOP_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0_CM8I,
      D3 => GRLFPC2_0_FPI_LDOP_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpAregLoadEn_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpAregLoadEn_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpBregLoadEn: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_FPI_LDOP_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3067,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpBregLoadEn_0: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_FPI_LDOP_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3067,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_RomxzSL2FromC: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SALSBs_0_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SALSBs_0_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SBLSBs_0_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SBLSBs_0_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3552,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SCLSBs_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS_CM8I(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN784_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_113_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SCLSBs_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SelInitRemBit: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_0_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_1_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_2_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_3_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_4_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_5_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlaregexp_ExpAregLC_1_1x: AND2A port map (
      A => GRLFPC2_0_FPI_LDOP_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlaregxz_un7_xzaregloaden: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(5),
      B => GRLFPC2_0_FPI_LDOP_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregexp_un6_expbregloaden: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregexp_un6_expbregloaden_0: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregxz_un5_xzbregloaden_1: OR3 port map (
      A => GRLFPC2_0_FPI_LDOP_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregxz_xzBregLC_1_2x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregxz_xzBregLC_1_0_2x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregxz_xzBregLC_1_0_0_2x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregxz_xzBregLC_1_0_1_2x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregxz_xzBregLC_1_1_2x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlcregxz_un8_inforcregsn: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN8_INFORCREGSN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(315),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(311),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(311),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(309),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(309),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(294),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(294),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(293),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(293),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(292),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(292),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(291),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(291),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(288),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(288),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(284),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(284),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(277),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(277),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(314),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3548);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(310),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3552);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(308),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3554);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(307),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3555);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(306),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3556);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(305),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3557);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(301),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3561);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(299),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3563);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(297),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3565);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(290),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3572);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(289),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3573);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(282),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3580);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(280),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(35),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(272),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(43),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3590);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(270),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(45),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3592);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(269),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(46),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3593);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(265),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(50),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3597);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3550_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3558_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3559_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(13),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3560_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(15),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3562_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3564_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3566_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(20),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3567_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(28),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3575_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3576_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3577_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3579_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(34),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3581_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(35),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3583_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(39),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3586_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(40),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3587_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3588_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3589_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(44),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3591_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3594_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(48),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3595_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3596_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3598_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3599_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3600_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3601_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3602_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3603_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(312),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(304),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(303),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(302),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(300),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(298),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(296),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(295),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(287),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(286),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(285),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(283),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(281),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(280),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(279),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(276),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(275),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(274),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(273),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(271),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(268),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(267),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(266),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(264),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(263),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(262),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(261),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(260),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_0_n_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(259),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_0_N_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_n_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N_CM8I(37),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_n_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N_CM8I(57),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_n_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(278),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_n_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(258),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_0: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_4: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_5: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_6: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_7: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_sn_m1_8: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(373),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(372),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_CM8I(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_2x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(371),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_6x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(367),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_9x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(364),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_10x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(363),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(362),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_12x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(361),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_13x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(360),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_14x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(359),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_15x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(358),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_16x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(357),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_17x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(356),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_18x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(355),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_19x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(354),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_20x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(353),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_21x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(352),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_22x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(351),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_23x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(350),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_24x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(349),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_25x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(348),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_26x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(347),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_27x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(346),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_28x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(345),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_29x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(344),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_30x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(343),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_31x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(342),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(341),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_33x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(340),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_34x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(339),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_35x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(338),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_36x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(337),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_37x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(336),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_38x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(335),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_39x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(334),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_40x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(333),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_41x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(332),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_42x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(331),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_43x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(330),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_44x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(329),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_45x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(328),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_46x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(327),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(326),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(325),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_49x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(324),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_50x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(323),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_51x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(322),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_52x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(321),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_53x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(320),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(319),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(318),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(317),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_n_9x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(364),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_n_10x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(363),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_n_26x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(347),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_n_50x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(323),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_117(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118(53),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_119(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_120(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_121(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(7),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_122(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_123(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_124(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_125(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_126(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_127(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_128(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_129(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_130(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_131(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_132(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_133(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_134(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_135(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_136(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_137(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_138(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_139(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_140(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_141(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_142(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_143(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_144(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_145(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_146(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_147(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_148(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_149(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_150(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_151(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_37x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(37),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_152(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_153(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_154(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_155(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_156(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_157(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_159(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_161(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_162(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_163(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_165(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_166(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_167(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_168(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(54),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(54),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_169(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_170(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_0(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_93(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN10_STKGEN_N,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_tz_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_TZ(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_2_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_TZ(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_2(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_4_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_STKOUT,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_2(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_4(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_5_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_4(57),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_14_142x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_QUOBITS(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_CM8I(142),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14(142));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_14_cm8i_142x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_CM8I(142));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_116(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_3,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_117(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(2),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_60x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118(53),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_61x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_119(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_119(52),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_62x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_120(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_120(51),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_63x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_121(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_121(50),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_64x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_122(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_122(49),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(64));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_65x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_123(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_123(48),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_66x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_124(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_124(47),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(66));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_67x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_125(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_125(46),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(67));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_68x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_126(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_126(45),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_69x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_127(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_127(44),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(69));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_70x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_128(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_128(43),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(70));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_71x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_129(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_129(42),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_72x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_130(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_130(41),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(72));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_73x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_131(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_131(40),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(73));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_74x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_132(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_132(39),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_75x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_133(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_133(38),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(75));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_76x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_134(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_134(37),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(76));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_77x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_135(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_135(36),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_78x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_136(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_136(35),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_79x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_137(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_137(34),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_80x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_138(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_138(33),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_81x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_139(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_139(32),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_82x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_140(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_140(31),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_83x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_141(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_141(30),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_84x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_142(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_142(29),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_85x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_143(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_143(28),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_86x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_144(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_144(27),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(86));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_87x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_145(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_145(26),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(87));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_88x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_146(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_146(25),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(88));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_89x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_147(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_147(24),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(89));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_90x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_148(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_148(23),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(90));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_91x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_149(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_149(22),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(91));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_92x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_150(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_150(21),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(92));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_93x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_151(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_151(20),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(93));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_94x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_152(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_0(37),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(94));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_95x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_153(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_153(18),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(95));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_96x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_154(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_154(17),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(96));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_97x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_155(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_155(16),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(97));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_98x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_156(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_156(15),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(98));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_99x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_157(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_157(14),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(99));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_100x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158(13),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(100));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_101x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_159(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_159(12),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(101));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_102x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160(11),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(102));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_103x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_161(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_161(10),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(103));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_104x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_162(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_162(9),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(104));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_105x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_163(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_163(8),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(105));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_106x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(106));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_107x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_165(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_165(6),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(107));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_108x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_166(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_166(5),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(108));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_109x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_167(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_167(4),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(109));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_110x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_168(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_168(3),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(110));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_111x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_169(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_169(2),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(111));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_112x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_170(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_170(1),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(112));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_113x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(113));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_49_258x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49(258));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_50_316x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_116(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_50(316));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_expybus_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_expybus_1_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_expybus_1_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0x: OR4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_1x: OR4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_CM8I(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_CM8I(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_4x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_6x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_7x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_10x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_11x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_12x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_14x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_15x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_16x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_17x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_19x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_21x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_22x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_23x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_24x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_26x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_29x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_30x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_35x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_37x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_39x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(39),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_42x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_43x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_44x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_45x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_46x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_47x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_48x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_49x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_50x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_51x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_53x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_55x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_57x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(55),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_n_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_N(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_2x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_3x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(8),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_10x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(10),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_11x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_12x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_14x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_15x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_16x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_17x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_19x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_21x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_22x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_23x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_24x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_26x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_29x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_30x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_35x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_37x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_39x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_42x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_43x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_44x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_45x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_46x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(42),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_47x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_48x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(44),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(48),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_49x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_50x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(46),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_51x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_53x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_55x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(55),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_56x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(56),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_57x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_10x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_11x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_12x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_14x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_15x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_16x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_17x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_19x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_21x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_22x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_23x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_24x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_26x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_29x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_30x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(25),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_35x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_37x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_39x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_42x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_43x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_44x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_45x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_46x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_47x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_48x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_49x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_50x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_51x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_53x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(55),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(55),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_56x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_57x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => N_5580,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232,
      S00 => N_5579,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => N_7993,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_CM8I(1),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_243,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_3x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3298,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3298,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(43),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SLCONTROL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_0_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_0_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_CM8I(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3295);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3298);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_2x: CM8 port map (
      D0 => N_7986,
      D1 => N_7986,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232,
      D3 => N_7986,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_245_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_269,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_0_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_d_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3295,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => N_5580);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_d_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S11 => NN_2,
      Y => N_7993);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_d_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S11 => NN_2,
      Y => N_7986);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_d_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_d_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_d_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_D_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_s_0x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_A7_0_N(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_CM8I(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_275,
      Y => N_5579);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_s_2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_2_CM8I(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_s_2_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_265,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_2_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_s_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_266,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_S_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_3_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_3_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_3_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_3_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_4_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_4_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_4_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_4_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_5_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_5_1x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_5_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_5_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_6_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_6(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_sn_m3_e: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(43),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN_N_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_gen_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(1),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN56_GEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_gen_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3548,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_gen_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_2: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2_CM8I,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_3: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3_CM8I,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un2_notprop: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(314),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(372),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un2_notprop_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3548,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un9_notprop_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(313),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un9_notprop_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(313),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un10_stkgen_n: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN10_STKGEN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un12_stkout: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un16_notprop: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3550_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un16_notprop_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un16_stkout: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_STKOUT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un22_gen: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN25_GEN,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un22_notprop: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un22_notprop_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un25_gen: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN392_CA_I,
      D1 => NN_4,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN392_CA_I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN25_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un28_notprop: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un28_notprop_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un35_notprop: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56(1),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un35_notprop_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un38_gen: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(1),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un38_gen_0: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56(1),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un42_notprop: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un47_gen: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN47_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un49_notprop: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un56_gen_0: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN56_GEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN784_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_113_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1_n_1x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N_CM8I(1),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN392_CA_I,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1_n_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3550_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_2_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_0_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_1_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_2_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_3_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_4_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_5_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_0_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_1_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_2_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_3_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_4_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_5_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_6_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_0_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_1_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_2_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_3_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_4_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_5_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_6: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_7: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_8: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_9: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_0: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_2: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_3: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_0: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_2: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_3: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_4: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_4_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_0: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_2: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_3: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_4: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_4_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_5: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_5_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notdivisorbit: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTDIVISORBIT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_4x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_6x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_7x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_7x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_1_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_0_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_1_0_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_2_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_2_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_2_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_2_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_2_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_3_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_3_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_3_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_3_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_3_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_4_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_4_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_4_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_4_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_5_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_5_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_5_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_5_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_6_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_6_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_6_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_6_8x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_7_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_7_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_7_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_8_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_8_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_8_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_9_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_9_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_9_6x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_10_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_10_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_11_4x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(0),
      S00 => GRLFPC2_0_FPO_FRAC(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(1),
      S00 => GRLFPC2_0_FPO_FRAC(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(2),
      S00 => GRLFPC2_0_FPO_FRAC_0(54),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_quobits_0x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_QUOBITS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_4x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(4),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(5),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_6x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(6),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_7x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(7),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(8),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_10x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(10),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_11x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_12x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(12),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(13),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_14x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(14),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_15x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(15),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_16x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(16),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_17x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(17),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(18),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_19x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(19),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(20),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_21x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(21),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_22x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(22),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_23x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(23),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_24x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(24),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(25),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_26x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(26),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(27),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(28),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_29x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(29),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_30x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(30),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(32),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(33),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(34),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_35x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(35),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(36),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_37x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(37),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(38),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(39),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_39x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(39),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(40),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(41),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_42x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(42),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_43x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(43),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_44x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(44),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_45x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(45),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_46x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(46),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_47x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(47),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(49),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(50),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(50),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(51),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(51),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(52),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(52),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(53),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(53),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(54),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(55),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(56),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(39),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_n_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N_CM8I(56),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N(57),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_n_57x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notsrres_1_n_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_0: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_3,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_0_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3288);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_2_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN54_SHDVAR_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN54_SHDVAR_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_2_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_STICKYFORSR1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_2_3: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN28_SHDVAR,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN10_SHDVAR,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_21x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_29x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_45x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_51x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(5),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_N(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_N(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I(57),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_N(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_n_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N_CM8I(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_n_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N_CM8I(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_n_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_n_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_n_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(244),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_n_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(242),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un10_shdvar: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(1),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN10_SHDVAR);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un24_shdvar_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un24_shdvar_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un24_shdvar_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1_CM8I,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un24_shdvar_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_STICKYFORSR1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un28_shdvar: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN28_SHDVAR);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un54_shdvar_1: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN54_SHDVAR_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un54_shdvar_4: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN54_SHDVAR_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectdivmult_un5_divmultv: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN5_DIVMULTV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectdivmult_un86_divmultv_n: OR4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTDIVISORBIT,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN86_DIVMULTV_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectdivmult_un111_divmultv: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTDIVISORBIT,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN111_DIVMULTV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectquobits_notdivc_1x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectquobits_notdivc_1_0x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_4_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4_CM8I(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4_CM8I(53),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_4_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_5_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5_CM8I(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5_CM8I(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_5_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_6_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6_CM8I(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(56),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(56),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6_CM8I(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3603_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_6_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_7_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7_CM8I(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7_CM8I(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3602_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_7_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_8_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8_CM8I(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(54),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(54),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8_CM8I(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3601_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_8_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_9_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9_CM8I(48),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9_CM8I(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3600_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_9_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_10_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10_CM8I(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10_CM8I(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3599_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_10_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_11_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11_CM8I(46),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11_CM8I(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3598_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_11_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_12_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12_CM8I(45),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_12_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3597,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_13_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13_CM8I(44),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13_CM8I(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3596_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_13_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_14_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14_CM8I(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14_CM8I(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3595_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_14_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_15_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15_CM8I(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15_CM8I(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3594_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_15_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_16_0_41x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_16_0_n_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0_N(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_17_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17_0(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17_CM8I(40),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_17_0_40x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17_0(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_17_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3592,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_18_0_39x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18_0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_19_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19_0(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19_CM8I(38),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_19_0_38x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19_0(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_19_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3590,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_20_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20_CM8I(37),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20_CM8I(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3589_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_20_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_21_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21_CM8I(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21_CM8I(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3588_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_21_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_22_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22_CM8I(35),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22_CM8I(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3587_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_22_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_23_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23_CM8I(34),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23_CM8I(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3586_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_23_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(39),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_24_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(38),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24_CM8I(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24_CM8I(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_24_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_25_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25_CM8I(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25_CM8I(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_25_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_26_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26_CM8I(31),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26_CM8I(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3583_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_26_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_27_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27_CM8I(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27_CM8I(30),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_27_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_28_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28_CM8I(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28_CM8I(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3581_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_28_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_29_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_0(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_CM8I(28),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_29_0_28x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_0(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_29_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3580,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_30_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30_CM8I(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30_CM8I(27),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3579_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_30_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_31_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(31),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31_CM8I(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31_CM8I(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_31_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_32_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32_CM8I(25),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32_CM8I(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3577_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_32_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_33_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33_CM8I(24),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33_CM8I(24),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3576_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_33_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_34_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34_CM8I(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34_CM8I(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3575_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_34_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_35_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35_CM8I(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35_CM8I(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(27),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_35_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_36_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(26),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(26),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36_CM8I(21),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_36_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3573,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_37_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37_0(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37_CM8I(20),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_37_0_20x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(25),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37_0(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_37_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3572,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_38_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(24),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38_CM8I(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(24),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_38_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_39_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39_CM8I(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39_CM8I(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_39_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_40_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(22),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40_CM8I(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(22),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_40_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_41_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(21),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41_CM8I(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41_CM8I(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(21),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_41_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_42_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42_CM8I(15),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42_CM8I(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3567_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_42_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_43_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43_CM8I(14),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43_CM8I(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3566_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_43_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_44_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_0(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_CM8I(13),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_44_0_13x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(18),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_44_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3565,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_45_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45_CM8I(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45_CM8I(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3564_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_45_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_46_11x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46_0(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46_CM8I(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_46_0_11x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(16),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_46_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3563,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_47_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47_CM8I(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47_CM8I(10),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3562_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_47_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_48_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48_0(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48_CM8I(9),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_48_0_9x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(14),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48_0(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_48_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3561,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_49_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49_CM8I(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49_CM8I(8),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3560_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_49_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_50_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50_CM8I(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50_CM8I(7),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3559_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_50_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_51_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51_CM8I(6),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51_CM8I(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3558_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_51_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_52_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(10),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52_CM8I(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_52_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3557,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_53_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_N(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53_CM8I(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_53_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3556,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_54_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_54_0_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_54_0_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(365),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_54_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_55_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_CM8I(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_55_0_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0_CM8I(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_55_0_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(366),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_55_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3554,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_56_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56_CM8I(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56_CM8I(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_56_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_61_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61_CM8I(52),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_61_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_62_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_CM8I(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_CM8I(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_3(54),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4(53),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_62_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_63_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63_CM8I(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_4(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_63_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_64_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64_CM8I(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64_CM8I(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_5(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_64_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_65_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65_CM8I(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65_CM8I(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_6(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_65_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_66_47x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66_0(47),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_7(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_66_0_47x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_67_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67_CM8I(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67_CM8I(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_8(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9(48),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_67_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_68_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68_CM8I(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68_CM8I(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_9(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10(47),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_68_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_69_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69_CM8I(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69_CM8I(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_69_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_70_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70_CM8I(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70_CM8I(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_11(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_70_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_71_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13(44),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71_CM8I(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71_CM8I(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_12(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_71_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_72_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72_CM8I(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72_CM8I(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_13(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_72_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_73_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73_CM8I(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73_CM8I(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_73_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_74_39x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0(39),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_74_0_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0_N(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16_0_N(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0_CM8I(39),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_74_0_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3593,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_75_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75_CM8I(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75_CM8I(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_16(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17(40),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_75_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_76_37x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0(37),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_76_0_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0_CM8I(37),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_3,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0_CM8I(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18_0(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3591_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_76_0_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_77_0_36x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19(38),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_77_0(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_78_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78_CM8I(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78_CM8I(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_19(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20(37),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_78_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_79_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79_CM8I(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79_CM8I(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_20(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_79_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_80_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80_CM8I(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80_CM8I(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_21(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22(35),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_80_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_81_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81_CM8I(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81_CM8I(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_22(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23(34),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_81_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_82_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_0(31),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_CM8I(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_0(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(37),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_82_0_31x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_82_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_0(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_83_30x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83_0(30),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_24(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_83_0_30x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83_0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_84_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84_CM8I(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84_CM8I(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN170_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_25_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_84_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_85_28x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85_CM8I(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ(30),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27(30),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_85_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_86_27x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86_CM8I(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ(29),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_86_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_87_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87_CM8I(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87_CM8I(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_28(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_87_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_88_0_25x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30(27),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88_0(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_89_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89_CM8I(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89_CM8I(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_30(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31(26),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_89_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_90_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90_CM8I(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90_CM8I(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_31(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32(25),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_90_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_92_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92_CM8I(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92_CM8I(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_33(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34(23),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_92_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_93_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93_CM8I(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93_CM8I(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_93_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_94_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94_CM8I(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_94_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_95_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95_CM8I(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95_CM8I(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_36(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37(20),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_95_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_96_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96_CM8I(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_37(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38(19),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_96_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_97_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97_CM8I(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97_CM8I(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_38(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39(18),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_97_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_98_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98_CM8I(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_39(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40(17),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_98_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_99_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99_CM8I(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99_CM8I(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_40(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41(16),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_99_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_100_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100_CM8I(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100_CM8I(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_41(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42(15),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_100_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_101_12x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101_CM8I(12),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ(14),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43(14),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_101_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_102_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102_CM8I(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102_CM8I(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_43(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_102_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_103_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103_CM8I(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103_CM8I(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_103_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_104_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104_CM8I(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104_CM8I(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_45(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_104_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_105_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105_CM8I(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105_CM8I(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47(10),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_105_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_106_7x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106_CM8I(7),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48(9),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_106_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_107_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107_CM8I(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107_CM8I(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_48(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_107_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_108_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108_CM8I(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108_CM8I(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_49(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_108_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_109_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109_CM8I(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109_CM8I(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_109_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_110_0_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_110_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_111_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111_CM8I(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_111_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_112_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112_CM8I(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_112_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_117_52x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_118_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_CM8I(51),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_118_0_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0_CM8I(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0_CM8I(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_118_0_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_118_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_119_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119_CM8I(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_61(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_119_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_119_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_120_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_CM8I(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_CM8I(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_62(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_120_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_121_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_CM8I(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_CM8I(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_63(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_121_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_122_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122_CM8I(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122_CM8I(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_64(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_122_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_123_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123_CM8I(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123_CM8I(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_65(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65(48),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_123_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_124_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124_CM8I(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124_CM8I(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_66(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66(47),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_124_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_125_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125_CM8I(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125_CM8I(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_67(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67(46),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_125_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_126_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126_CM8I(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126_CM8I(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_68(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_126_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_127_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127_CM8I(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127_CM8I(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_69(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_127_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_128_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128_CM8I(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128_CM8I(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_70(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_128_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_129_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_CM8I(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_CM8I(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_71(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_129_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_130_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_CM8I(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_CM8I(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_72(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72(41),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_130_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_131_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131_CM8I(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131_CM8I(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_73(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73(40),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_131_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_132_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132_CM8I(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132_CM8I(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_74(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_132_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_133_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133_CM8I(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133_CM8I(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_75(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_133_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_134_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134_CM8I(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134_CM8I(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_76(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76(37),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_134_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_135_34x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0(34),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_77(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_135_0_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0_CM8I(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0_CM8I(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_77_0(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_18(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_135_0_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_136_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136_CM8I(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136_CM8I(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_78(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78(35),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_136_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_137_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_CM8I(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_CM8I(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_79(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79(34),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_137_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_138_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138_CM8I(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138_CM8I(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_80(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_138_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_139_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139_CM8I(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139_CM8I(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81(32),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_139_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_140_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_CM8I(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_CM8I(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_82(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_140_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_141_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141_CM8I(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141_CM8I(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN574_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83_0(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_141_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_142_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142_CM8I(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142_CM8I(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84(29),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_142_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_143_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143_CM8I(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143_CM8I(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_143_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_144_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144_CM8I(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144_CM8I(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_86(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86(27),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_144_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_145_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145_CM8I(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145_CM8I(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_87(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87(26),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_145_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_146_23x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0(23),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_88(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_146_0_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0_CM8I(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0_CM8I(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88_0(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_29(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_146_0_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_147_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147_CM8I(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147_CM8I(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_89(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89(24),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_147_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_148_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148_CM8I(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148_CM8I(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_148_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_149_20x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0(20),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_91(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_149_0_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0_CM8I(20),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0_CM8I(20),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N(24),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_149_0_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_150_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_CM8I(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_92(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_150_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_151_0_18x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93(20),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_0(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_152_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152_CM8I(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_94(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94(19),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_152_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_153_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153_CM8I(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153_CM8I(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_95(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95(18),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_153_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_154_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_CM8I(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_96(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96(17),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_154_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_155_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155_CM8I(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155_CM8I(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_97(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97(16),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_155_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_156_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156_CM8I(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156_CM8I(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_98(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98(15),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_156_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_157_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157_CM8I(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157_CM8I(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_99(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99(14),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_157_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_158_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_CM8I(11),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43(14),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ(14),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_0(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_158_0_11x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100(13),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_158_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_159_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159_CM8I(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159_CM8I(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_101(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_159_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_160_9x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160_CM8I(9),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_160_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_161_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161_CM8I(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161_CM8I(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_103(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_161_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_162_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162_CM8I(7),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162_CM8I(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_104(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104(9),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_162_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_163_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163_CM8I(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163_CM8I(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105(8),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_163_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_164_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164_CM8I(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_164_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_165_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165_CM8I(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165_CM8I(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_107(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_165_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_166_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166_CM8I(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166_CM8I(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_108(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_166_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_167_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167_CM8I(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_109(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_167_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_168_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_110(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_168_0_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0_CM8I(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_110_0(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_168_0_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SALSBs_1_0_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0_CM8I(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SALSBs_1_0_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(369),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SBLSBs_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_CM8I(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SBLSBs_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SCLSBs_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1_CM8I(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_112_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SCLSBs_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN681_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN678_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N_CM8I,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN165_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN507_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN339_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN336_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN336_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN339_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_un339_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN339_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_un392_ca_i: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN392_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_un681_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_UN681_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_CA_56_1x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SALSBS_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_56(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_CA_113_0_1x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_56(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_113_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_CA_170_1x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_112(1),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_112_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_CA_170(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN678_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN675_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN336_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN333_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN333_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN336_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN507_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN504_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN504_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN507_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN165_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN162_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un165_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN165_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un336_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN336_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un507_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN507_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un678_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN678_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un784_ca_i: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_UN784_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_55_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3552,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55_CM8I(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55_CM8I(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_55_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_55_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_112_0_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_54(3),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_112_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_169_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_111(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_111(3),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_CA_169(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN675_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN672_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN333_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN330_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN330_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN333_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN504_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN162_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un162_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN162_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un333_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN333_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un504_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN504_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un675_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN675_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un777_ca_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I_CM8I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un777_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_UN777_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_CA_54_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_54(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_CA_111_3x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53(4),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_111(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_CA_168_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_110(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_0(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_168(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN672_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN669_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N_CM8I,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_CIN_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN498_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN498_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN330_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN156_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_un330_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN330_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_un672_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_UN672_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_53_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3554,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53_CM8I(4),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53_CM8I(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_53_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_53_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_110_4x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52(5),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_110(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_167_4x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_109(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_109(5),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_CA_167(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_0_1(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN156_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN498_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN495_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN495_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN498_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN669_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN666_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN324_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un156_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN156_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un498_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN498_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un669_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_UN669_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_52_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3555,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52_CM8I(5),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52_CM8I(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_52_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_54_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_52_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_109_5x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51(6),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_52(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_109(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_166_5x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_108(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_108(6),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108(5),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_CA_166(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN666_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN663_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN495_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN492_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN150_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN324_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN321_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN321_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN324_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un324_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN324_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un495_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN495_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un666_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_UN666_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_51_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(9),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51_CM8I(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_51_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3556,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_51_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_108_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50(7),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50(7),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_108(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_165_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_107(7),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_107(7),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_CA_165(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN663_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN660_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN492_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN489_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN150_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN321_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un150_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN150_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un321_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN321_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un492_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN492_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un663_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_UN663_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_50_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(10),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(10),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50_CM8I(7),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_50_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3557,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_50_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_107_7x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_49(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_49(8),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_107(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_164_0_7x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_164_0_tz_7x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_48(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ_CM8I(7),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_164_0_tz_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_CA_164_0_TZ_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN489_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN486_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN144_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN660_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN657_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN315_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un489_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN489_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un660_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN660_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un1141_ca_i: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_CIN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_48(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un1141_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_UN1141_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_CA_49_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(11),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(11),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3558_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_49(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_CA_163_8x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105(9),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_CA_163(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN657_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN654_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_0(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN486_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN483_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN144_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN315_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un144_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN144_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un315_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN315_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un486_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN486_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un657_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_UN657_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_48_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(12),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3559_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_48(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_105_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48(9),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_105_0_tz_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_3,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ_CM8I(9),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(13),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_105_0_tz_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_105_0_TZ_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_162_9x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_104(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_104(10),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_CA_162(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN654_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN651_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN138_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN138_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN483_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN480_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN480_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN483_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN309_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un483_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN483_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un654_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN654_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un728_ca_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un728_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_UN728_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_CA_104_10x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46(11),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_104(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_CA_161_10x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_103(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_103(11),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_CA_161(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN138_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN309_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN480_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN477_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN477_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN480_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN651_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN648_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un138_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN138_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un309_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN309_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un480_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN480_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un651_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_UN651_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_46_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(14),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46_CM8I(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_46_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3561,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_46_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_103_11x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_45(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_45(12),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_103(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_160_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_160_0_tz_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44(13),
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ_CM8I(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_160_0_tz_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_CA_160_0_TZ_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN648_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN645_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN477_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN474_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN132_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN303_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN303_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un477_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN477_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un648_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN648_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un1113_ca_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44(13),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un1113_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_UN1113_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_CA_45_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(15),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3562_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_45(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_CA_159_12x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_101(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_101(13),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_CA_159(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN645_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN642_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN474_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN471_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN303_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN300_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN132_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un132_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN132_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un303_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN303_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un474_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN474_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un645_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN645_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_44_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(16),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(16),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44_CM8I(13),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_44_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3563,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_44_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_101_13x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_43(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_43(14),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_101(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_158_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158_CM8I(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158_0(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_158_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_CA_158_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN300_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN297_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN471_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN468_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN642_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN639_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN126_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un300_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN300_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un471_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN471_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un642_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN642_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_43_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3564_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_43(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_100_0_tz_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(18),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ_CM8I(14),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_0(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_100_0_tz_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_100_0_TZ_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_157_14x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_99(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_99(15),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_CA_157(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN468_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN465_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN639_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN636_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN126_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN123_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN297_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN294_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un126_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN126_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un297_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN297_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un468_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN468_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un639_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN639_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un693_ca_i: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(18),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44_0(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un693_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN693_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_CA_99_15x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_41(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_41(16),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_99(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_CA_156_15x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_98(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_98(16),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_CA_156(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN636_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN633_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN294_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN291_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN123_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN120_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN465_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN462_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un123_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN123_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un294_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN294_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un465_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN465_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un636_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN636_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_CA_41_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(19),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3566_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_41(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_CA_98_16x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_40(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_40(17),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_98(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_CA_155_16x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_97(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_97(17),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_CA_155(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN291_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN288_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN462_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN459_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN633_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN630_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN120_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un120_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN120_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un291_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN291_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un462_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN462_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un633_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN633_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_CA_40_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(20),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(20),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3567_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_40(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_CA_97_17x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_39(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_39(18),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_97(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_CA_154_17x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_96(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_96(18),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_96(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_CA_154(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN459_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN456_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN288_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN285_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN630_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN627_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_1(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN114_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN114_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un288_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN288_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un459_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN459_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un630_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_UN630_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_CA_39_18x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(21),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_39(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_CA_96_18x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_38(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_38(19),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_96(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_CA_153_18x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_95(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_95(19),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_CA_153(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN627_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN624_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN285_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN282_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN114_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN111_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN456_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN453_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_un114_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN114_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_un285_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN285_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_un456_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN456_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_un627_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_2(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_UN627_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_CA_38_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_38(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_CA_95_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_37(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_37(20),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_38(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_95(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_CA_152_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_94(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_94(20),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_CA_152(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN453_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN450_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN282_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN279_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN111_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN108_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN624_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN621_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_un111_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN111_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_un282_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN282_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_un453_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN453_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_un624_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_UN624_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_CA_37_20x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(23),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_37(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_CA_94_20x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_36(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_36(21),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_94(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_CA_151_20x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_93(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_93(21),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_93(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_CA_151(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN621_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN618_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN450_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN447_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN108_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN105_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN279_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un108_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN108_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un279_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN279_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un450_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN450_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un621_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_UN621_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_CA_36_21x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(24),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_36(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_CA_93_21x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35(22),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_93(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_CA_150_21x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_92(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_92(22),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_92(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_CA_150(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN618_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN615_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN447_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN444_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN105_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN273_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un105_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN105_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un447_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN447_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un618_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_UN618_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_35_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(25),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35_CM8I(22),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_6,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_35_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3572,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_35_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_92_22x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34(23),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_35(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_92(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_149_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_91(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_0(20),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_CA_149(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN444_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN441_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN615_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN612_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN99_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN273_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN270_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN270_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN273_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un273_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN273_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un444_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN444_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un615_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_UN615_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_34_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34_CM8I(23),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_34_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3573,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_34_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_91_23x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_33(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_33(24),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_91(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_148_23x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_CA_148(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN270_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN267_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN612_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN609_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN441_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN99_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un99_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN99_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un270_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN270_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un441_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN441_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un612_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_UN612_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_33_24x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(27),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_33(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_90_0_24x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N(24),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_33(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_90_0_tz_n_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34(23),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N_CM8I(24),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(28),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_90_0_tz_n_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_90_0_TZ_N_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_147_24x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_89(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_89(25),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_CA_147(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN267_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN264_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_3(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN609_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN606_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN93_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN93_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN435_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un267_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN267_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un609_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN609_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un623_ca_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_34(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un623_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_UN623_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_CA_89_25x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_31(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_31(26),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_89(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_CA_146_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_88(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146_0(23),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_CA_146(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN606_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN603_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN264_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN261_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN435_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN432_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_3_n: OR2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_CIN_3_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN93_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN90_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un93_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN93_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un264_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN264_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un435_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN435_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un606_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_UN606_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_CA_31_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(29),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3576_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_31(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_CA_88_26x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_30(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_30(27),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_88(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_CA_145_26x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_87(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_87(27),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_CA_145(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN261_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN258_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN432_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN429_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN603_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN600_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_2(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN90_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN87_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un90_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN90_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un261_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN261_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un432_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN432_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un603_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_UN603_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_CA_30_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(30),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(30),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3577_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_30(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_CA_87_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_30(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_29(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88_0(25),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_87(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_CA_144_27x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_86(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_86(28),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_CA_144(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN429_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN426_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN600_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN597_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN258_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN255_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN87_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN84_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un87_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN87_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un258_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN258_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un429_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN429_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un600_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_UN600_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_CA_29_28x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(31),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_29(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_CA_86_28x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_28(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_28(29),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_86(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_CA_143_28x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85(29),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_CA_143(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN597_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN594_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN84_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN81_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN426_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN423_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN255_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN252_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un84_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN84_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un255_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN255_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un426_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN426_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un597_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_UN597_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_28_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3579_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_28(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_85_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_85_0_tz_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(33),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ_CM8I(29),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_0(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_85_0_tz_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_85_0_TZ_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_142_29x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84(30),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_CA_142(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN594_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN591_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN423_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN420_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN81_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN78_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_7,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN252_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN249_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un81_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN81_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un252_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN252_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un423_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN423_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un588_ca_i: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(33),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29_0(28),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un588_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN588_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un594_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_UN594_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_84_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27(30),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_84_0_tz_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_1,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ_CM8I(30),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(34),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_84_0_tz_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_84_0_TZ_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_141_30x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83(31),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_CA_141(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN591_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN588_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN249_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN246_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN78_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN420_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN417_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un78_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN78_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un249_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN249_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un420_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN420_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un581_ca_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(34),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un581_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_CIN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN581_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un591_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_UN591_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_CA_83_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN170_CA_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_25_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_CA_83_0_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_25_0(32),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN170_CA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_83_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_CA_140_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_82(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_82(32),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_CA_140(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN588_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN585_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN246_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN243_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN72_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN417_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un246_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN246_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un417_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN417_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un574_ca_i: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_25_0(32),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN170_CA_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN574_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un588_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_UN588_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_CA_25_0_32x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_25_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_CA_82_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_24(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83_0(30),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_82(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_CA_139_32x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81(33),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_CA_139(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN585_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN582_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN243_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN411_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_3(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN72_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_3(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un72_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN72_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un170_ca_i: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3582,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN170_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un243_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN243_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un585_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_UN585_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_24_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3583_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_24(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_81_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_24(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81_CM8I(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82_0(31),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_81_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_82(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_81_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_138_33x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_80(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_80(34),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_CA_138(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN582_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN579_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN411_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN408_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN66_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN66_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN237_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN237_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_4(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_un411_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN411_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_un582_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_UN582_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_CA_80_34x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_22(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_22(35),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_80(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_CA_137_34x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_79(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_79(35),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_79(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_CA_137(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN579_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN576_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN66_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN63_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN408_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN405_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN237_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN234_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un66_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN66_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un237_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN237_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un408_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN408_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un579_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_UN579_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_CA_22_35x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_22(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_CA_79_35x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_21(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_21(36),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_79(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_CA_136_35x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_78(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_78(36),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_CA_136(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN234_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN231_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN576_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN573_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN405_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN402_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN63_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un63_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN63_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un234_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN234_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un405_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN405_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un576_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_UN576_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_CA_21_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(39),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3586_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_21(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_CA_78_36x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_20(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_20(37),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_21(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_78(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_CA_135_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_77(37),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_0(34),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_CA_135(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN231_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN228_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN402_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN399_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN573_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN570_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN57_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un231_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN231_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un402_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN402_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un573_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_4(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_UN573_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_CA_20_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3587_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_20(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_CA_77_37x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_19(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_19(38),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_77(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_CA_134_37x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_76(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_76(38),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_CA_134(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN228_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN225_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN570_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN567_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN57_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN399_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN396_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un57_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN57_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un228_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN228_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un399_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN399_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un570_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_UN570_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_CA_19_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(41),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3588_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_19(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_CA_76_38x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_18(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_18(39),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_19(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_76(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_CA_133_38x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_75(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_75(39),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_CA_133(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_cin_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN567_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN564_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN51_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN225_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN222_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN396_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_un225_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN225_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_un396_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_7(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN396_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_un567_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_UN567_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_CA_18_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3589_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_18(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_CA_75_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17(40),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76_0(37),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_75(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_CA_132_39x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_74(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_74(40),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_CA_132(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_cin: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN564_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN561_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN222_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN219_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN51_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN48_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN390_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_un51_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN51_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_un222_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN222_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_un564_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_UN564_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_17_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(43),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17_CM8I(40),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_17_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3590,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_17_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_74_40x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_16(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_16(41),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_74(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_131_40x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_73(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_73(41),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_CA_131(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN219_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN216_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN561_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN558_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN390_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN387_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN48_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un48_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN48_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un219_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN219_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un390_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN390_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un561_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_UN561_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_CA_16_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(44),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3591_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_16(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_CA_73_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15(42),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74_0(39),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_73(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_CA_130_41x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_72(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_72(42),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_72(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_CA_130(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN216_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN213_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN558_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN555_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN387_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN384_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN42_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN42_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_4(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un216_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN216_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un387_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN387_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un558_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_UN558_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_15_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(45),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15_CM8I(42),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_15_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3592,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_15_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_72_42x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14(43),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_72(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_129_42x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_71(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_71(43),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_71(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_CA_129(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN384_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN381_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN555_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN552_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN42_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN39_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN213_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN210_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_5(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un42_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN42_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un213_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN213_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un384_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN384_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un555_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_UN555_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_14_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(46),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14_CM8I(43),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_14_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3593,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_14_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_71_43x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_13(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_13(44),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_14(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_71(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_128_43x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_70(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_70(44),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_CA_128(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN381_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN378_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN39_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN39_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN210_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN207_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN552_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN549_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un39_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN39_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un210_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN210_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un381_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN381_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un552_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_UN552_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_CA_13_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(47),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3594_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_13(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_CA_70_44x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_12(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_12(45),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_13(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_70(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_CA_127_44x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_69(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_69(45),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_CA_127(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN549_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN546_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_4(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN378_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN375_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN33_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN33_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN207_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN204_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN204_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN207_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_3(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un207_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN207_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un378_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN378_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un549_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_UN549_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_CA_12_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(48),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3595_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_12(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_CA_69_45x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_11(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_11(46),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_69(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_CA_126_45x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_68(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_68(46),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_CA_126(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN375_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN372_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN546_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN543_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN33_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN30_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN204_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN201_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN201_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN204_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un33_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN33_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un204_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN204_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un375_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN375_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un546_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_5(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_UN546_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_CA_11_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(49),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3596_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2_8,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_11(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_CA_68_46x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10(47),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_68(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_CA_125_46x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_67(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_67(47),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_CA_125(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN372_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN369_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN543_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN540_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN30_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN27_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN201_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN198_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN198_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN201_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un30_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN30_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un201_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN201_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un372_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN372_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un543_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_UN543_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_10_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(50),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10_CM8I(47),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_10_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3597,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_10_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_67_47x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_9(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_9(48),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_10(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_67(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_124_47x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_66(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_66(48),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_CA_124(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN369_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN366_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN540_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN537_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN198_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN27_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN24_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un27_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN27_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un198_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN198_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un369_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_8(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN369_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un540_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_UN540_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_CA_9_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(51),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3598_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_9(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_CA_66_48x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_8(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_8(49),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_66(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_CA_123_48x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_65(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_65(49),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_CA_123(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN366_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN363_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN192_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN192_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN24_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN21_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN537_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN534_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_un24_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN24_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_un366_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN366_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_un537_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_UN537_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_CA_8_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(52),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3599_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_CA_65_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_7(50),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66_0(47),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_65(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_CA_122_49x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_64(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_64(50),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_CA_122(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN363_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN360_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN534_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN531_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN21_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN192_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN189_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_un21_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN21_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_un192_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN192_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_un363_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN363_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_un534_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_UN534_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_CA_7_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(53),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(53),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3600_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_7(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_CA_64_50x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_6(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_6(51),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_64(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_CA_121_50x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_63(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_63(51),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_CA_121(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN189_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN186_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_6(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN531_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN528_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_cin_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO_4,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN15_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN360_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN357_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_5(2),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un189_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN189_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un360_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN360_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un531_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_UN531_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_CA_6_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(54),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3601_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_6(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_CA_63_51x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_5(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_5(52),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_63(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_CA_120_51x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_62(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_62(52),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_CA_120(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN357_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN354_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN186_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN183_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN528_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN525_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN15_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN12_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un15_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN15_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un186_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN186_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un357_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN357_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un528_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_UN528_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_CA_5_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3602_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_5(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_CA_62_52x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_4(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_4(53),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_5(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_62(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_CA_119_52x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_61(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_61(53),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_61(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_CA_119(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN183_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN180_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN354_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN351_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN12_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN525_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN522_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un12_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN12_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un183_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN183_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un354_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN354_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un525_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_UN525_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_4_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(56),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(56),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3603_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_SN_N_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_4(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_61_53x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_3(54),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_3(54),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_61(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_118_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118_CM8I(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118_0(51),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_118_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_118(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_CA_118_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN180_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN177_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN351_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN348_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN6_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN6_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_10(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN522_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN519_TEMP,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT_5(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un180_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN180_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un351_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN351_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un522_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_UN522_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_3_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_3(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_60_0_tz_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ_CM8I(54),
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4(53),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_60_0_tz_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_117_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_59(55),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_59(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_117(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN519_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN516_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN177_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN6_TEMP,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN348_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN345_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN345_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN348_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_11(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un6_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN6_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un177_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN177_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un348_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN348_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un519_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_6(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_UN519_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_CA_59_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_CA_60_0_TZ(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_59(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_CA_116_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_59(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_116(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN516_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN513_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN79_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_temp2_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN171_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_temp2_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN345_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN342_TEMP,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN342_TEMP,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN345_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un345_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_9(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN345_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un408_ca_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un408_ca_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN408_CA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un516_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_UN516_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_cin_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_cin_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN171_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN171_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(3),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN513_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un171_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP_1_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN171_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un228_sa_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4_N(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_4(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un228_sa_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un342_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN342_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un456_sa_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN31_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_59(55),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un456_sa_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN228_SA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un513_temp: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTMULTIP(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN513_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un684_sa_i: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN55_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_CA_116(55),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un684_sa_i_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN456_SA_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_UN684_SA_I_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_CM8I(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_3,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_111(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_57_0_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN8_ZERO,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_57_0_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(368),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_57_0_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_113_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_CM8I(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_CA_54(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_55(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_113_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_CIN_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_CM8I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_6: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_7: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_0: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_1: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_3: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_4: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_5: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden_0: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden_1: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden_2: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden_3: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden_4: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden_5: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_entrypoint_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN5_S_0,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1500,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0_CM8I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_entrypoint_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_s_cmp_1: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_s_cmp_1_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_entrypoint: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_14_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_0_N,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_0_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_entrypoint_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_s_14_0_n: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4260,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_0_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_s_dyadic_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un5_s_0: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN5_S_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un9_s_14_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_14_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un14_s_mov_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_computeconst_un49_resvec: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      B => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_1_6x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3678);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_1_9x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3681);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_CM8I(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_1x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_3x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_EXPYBUS_1(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_4x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_5x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3678,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3678,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_7x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3681,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_8x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3681,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_9x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3681,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_10x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_11x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_12x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expybus_2_2x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_mixoin_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(35),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_0x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_1x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_2x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_3x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_4x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3713,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_5x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3714,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_6x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3715,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_7x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3716,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_8x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3717,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_9x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3718,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_10x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I(10),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_11x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I(11),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_12x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I(12),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un40_expxbus_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3275_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_0_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3286,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3286,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3279,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3278,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_6_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_6_N_CM8I,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_6_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_6_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_6_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_7_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7_N_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3282,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_6_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_7_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_9: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3277,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_9_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_stickyforsr1: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_STICKYFORSR1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_NOTXZYFROMD,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_NOTXZYFROMD,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un5_notxzyfromd: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_NOTXZYFROMD);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un5_xzybuslsbs: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(1),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(1),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3378,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3434_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_3x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(3),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_4x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_5x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_6x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3383,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3439_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_8x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_9x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(9),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3386,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3442_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3387,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3443_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_12x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(12),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_13x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(13),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_14x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(14),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3391,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3447_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_16x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(16),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_17x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_18x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(18),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_19x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(19),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3396,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3452_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_21x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(21),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_22x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(22),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_23x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(23),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_24x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(24),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_25x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(25),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_26x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(26),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3403,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3459_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_28x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(28),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_29x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(29),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3406,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3462_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_31x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(31),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_32x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(32),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_33x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(33),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_34x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(34),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3411,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3467_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3412,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3468_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3413,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3469_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_38x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(38),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_39x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(39),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_40x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(40),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_41x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(41),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_42x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3419,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3475_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_44x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(44),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_45x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(45),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3422,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3478_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_47x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(47),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_48x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(48),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3425,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3481_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3426,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3482_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_51x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(51),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3428,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3484_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_53x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(53),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_54x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(54),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_55x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(55),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_56x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(56),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(57),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3489_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un19_xzxbus_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN26_NOTXZYFROMD,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_6: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_7: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_8: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_9: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_10: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_11: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_12: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un26_notxzyfromd: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN26_NOTXZYFROMD);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un37_notxzyfromd: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un37_notxzyfromd_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_55,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_2: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(57),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3310_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(57),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3365_I_0,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3365_I_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(56),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(56),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_5: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3314_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_7: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(31),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3322_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_9: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(26),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3335_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_11: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3338_I_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_7,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(29),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_11_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1812_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_12: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3313_I_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(13),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_12_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1796_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_13: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13_CM8I,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3316_I_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(44),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_13_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_15_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3347,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3347,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_17: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(51),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_17_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3319,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_19: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(54),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(54),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_19_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3324,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_24: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_24_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_25: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_25_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3342,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_28: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(34),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_28_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3333,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_29: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29_CM8I,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_29_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3331,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_31_n: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3327,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3327,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_34: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(27),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_34);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_36: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3340,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3312,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3334_I_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_9,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_37: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3326,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_37_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_39: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(35),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3355_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(35),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_39_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_41: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(43),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3357_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_41_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_42: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(10),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42_S,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_42_s: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42_S_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3350,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3351,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42_S);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_42_s_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_1831_S,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42_S_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_43: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3363_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_43_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_45: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3346,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_45_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_46: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3360,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_48: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3318,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3325,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_48);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_50_n: OR4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3348,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3356,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_51: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3329,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3330,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_55: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_34,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_55);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_56: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_48,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_56_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_1x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_32x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_33x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_34x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_35x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_37x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_38x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_39x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_40x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_41x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_42x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_43x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_44x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_45x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_46x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_47x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_49x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_50x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_51x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_52x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_53x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_54x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2_30x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2_0_30x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2_1_30x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2_2_30x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3379,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3380,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3381,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3382,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3384,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3385,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(9),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3388,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(12),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3389,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(13),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3390,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(14),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3392,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(16),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3393,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(17),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3394,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(18),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3395,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3397,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(21),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3398,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(22),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3399,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(23),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3400,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(24),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3401,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(25),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3402,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(26),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3404,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(28),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3405,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(29),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3407,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3408,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(32),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3409,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(33),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3410,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(34),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3414,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(38),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3415,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(39),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3416,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(40),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3417,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(41),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3418,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(42),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3420,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(44),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3421,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(45),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3423,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(47),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3424,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3427,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(51),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3429,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(53),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3430,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(54),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3431,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(55),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3432,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(56),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3378);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3379);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3380);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3381);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3382);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3383);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3384);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3385);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3386);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3387);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3388);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3389);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3390);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3391);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3392);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3393);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3394);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3395);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3396);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3397);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3398);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3399);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3400);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3401);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_7,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3402);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3403);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3404);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3405);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3406);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3407);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3408);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3409);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3410);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_8,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3411);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3412);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3413);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3414);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3415);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3416);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3417);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3418);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3419);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_9,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3420);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3421);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3422);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3423);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3424);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3425);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3426);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3427);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3428);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_10,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3429);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3430);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3431);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_0_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3432);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_2x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(229),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3434_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_7x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(224),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3439_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_10x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(221),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3442_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_11x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(220),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3443_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_15x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(216),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3447_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_20x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(211),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_11,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3452_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_27x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(204),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3459_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_30x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(201),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3462_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_35x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(196),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3467_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_36x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(195),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3468_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_37x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(194),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3469_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_43x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(188),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3475_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_46x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(185),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3478_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_49x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(182),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3481_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_50x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(181),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_12,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3482_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_52x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(179),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3484_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_1_n_57x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(174),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3489_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(15),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_STICKYFORSR1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_CM8I(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(231),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(230),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(228),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(227),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(226),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(225),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(223),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(222),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(219),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(218),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(217),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(215),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(214),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(213),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(212),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(210),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(209),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(208),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(207),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(206),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(205),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(203),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(202),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(200),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(199),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(198),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(197),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(193),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(192),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(191),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(190),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(189),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(187),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(186),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(184),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(183),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(180),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(178),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(177),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(176),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(175),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0_1: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0_2: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0_3: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0_4: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m2_0_5: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M2_0_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_0_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_0_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_1_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_1_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_2_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_2_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_2_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_2_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_3_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_3_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_3_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_3_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_4: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_4_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_4_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_4_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_4_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_5: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_5_CM8I,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_5_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3490_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_5_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_5_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m4_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN37_NOTXZYFROMD,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_M4_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_notam2_0: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un2_inexact: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_CM8I,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un2_inexact_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STATUS_1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un2_inexact_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un13_inexact_0_n: OR2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STATUS_1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_0_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_0: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_1: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_2: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_3: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_4: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_5: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_10: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_11: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_15: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_15_CM8I,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_15_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_15_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_16: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_16_CM8I,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_16);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_16_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_16_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_21: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_21);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_22_n: OR3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_22_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_25: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_11,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_25_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_10,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_25_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_25_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_26: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_21,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_16,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_15,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_26);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_27: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_27_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_22_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_27);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_27_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_27_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notabortnullexc: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_TEMP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_4_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_4_0_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_4_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2662);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_4_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_4_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_6_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2662,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_6_0_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2664);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_6_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_6_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_7_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_7_0_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2664,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2664,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2665);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_7_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_7_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_10_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_10_0_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(244),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2668);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_10_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_10_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_13_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_13_0_CM8I,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_13_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2671);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_13_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_13_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_15_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2665,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2668,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2671,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2673);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_17_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2675);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_20_0: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2678);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_21_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_21_0_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2678,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2678,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2679);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_21_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_21_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_23_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_23_0_CM8I,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_23_0_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_23_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(9),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(7),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN4_LOCUV,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2681);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_23_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_23_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_d: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_0_D_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      D2 => N_7976,
      D3 => N_7976,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1,
      S01 => NN_4,
      S10 => N_5581,
      S11 => N_7971_N,
      Y => N_7974);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_d_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_0_D_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_d_d_1: CM8 port map (
      D0 => N_8050,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2673,
      D2 => N_8050,
      D3 => N_8050,
      S00 => N_7971_N,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      S11 => N_5577,
      Y => N_7976);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_d_d_1_d_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2675,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2679,
      S00 => N_7971_N,
      S01 => NN_4,
      S10 => N_5577,
      S11 => NN_2,
      Y => N_8050);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_s: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      Y => N_5577);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_s_0: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      Y => N_5581);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_s_2_n: CM8 port map (
      D0 => N_5577,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      S00 => N_5581,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_0_S_2_N_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      Y => N_7971_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_s_2_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_0_S_2_N_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_27_0_s_3: AND2 port map (
      A => N_5581,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      Y => N_7973);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0: CM8 port map (
      D0 => N_7974,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2681,
      D2 => NN_4,
      D3 => NN_4,
      S00 => N_7973,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_0: CM8 port map (
      D0 => N_7974,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2681,
      D2 => NN_4,
      D3 => NN_4,
      S00 => N_7973,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_oprexcshft_un3_oprexc: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_6(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_N,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(58),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_CM8I(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(58),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      S11 => GRLFPC2_0_FPO_FRAC_0(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(57),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_n_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_N_CM8I(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_N(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_n_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_N_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_u_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(59),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN4_LOCUV,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedbackmulxff_un18_feedback: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedbackmulxff_un19_feedback: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_mapmulxff_unimpmap: CM8 port map (
      D0 => cpi_d_inst(13),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP_CM8I,
      D2 => NN_4,
      D3 => cpi_d_inst(12),
      S00 => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
      S01 => cpi_d_inst(9),
      S10 => cpi_d_inst(19),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_mapmulxff_unimpmap_cm8i: CM8INV port map (
      A => cpi_d_inst(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_exmiptr_2x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_EXMIPTR(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_0_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(1),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2025);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_0_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_0_n_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_N,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK_N(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0(3),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_0_N_CM8I(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2024_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_0_n_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_0_N_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(1),
      D1 => cpi_d_inst(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2034);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(2),
      D1 => cpi_d_inst(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2035);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(3),
      D1 => cpi_d_inst(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2036);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(4),
      D1 => CPI_D_INST_0(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2037);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(5),
      D1 => cpi_d_inst(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2038);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(6),
      D1 => cpi_d_inst(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2039);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(7),
      D1 => cpi_d_inst(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2040);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_1_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(8),
      D1 => cpi_d_inst(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2041);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2036,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_EXMIPTR(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2046);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2037,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2037,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2047);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2038,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2048);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2039,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2049);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2041,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(7),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2051);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_2_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_sn_m2_0_a2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN4_TEMP2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_sn_m2_0_a2_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN4_TEMP2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_sn_m4_i: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_SN_N_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_sn_m6_0_a2: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN4_NOTRESETORUNIMP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_sn_m6_0_a2_0: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN4_NOTRESETORUNIMP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_pctrl_new_2_0_65x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(64),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_2_0(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_pctrl_new_14_77x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_2(77),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_pctrl_new_14_0_77x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_2(77),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_0(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_pctrl_new_14_2_77x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(46),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_TEMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_2(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_un4_temp2: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(63),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN4_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un4_locuv: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN4_LOCUV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un20_locov_3_n: OR3C port map (
      A => GRLFPC2_0_FPO_EXP(2),
      B => GRLFPC2_0_FPO_EXP(1),
      C => GRLFPC2_0_FPO_EXP(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_3_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un20_locov_5: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_FPO_EXP(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_FPO_EXP(6),
      S01 => GRLFPC2_0_FPO_EXP(5),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_3_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un20_locov_5_cm8i: CM8INV port map (
      A => GRLFPC2_0_FPO_EXP(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un21_locov: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_FPO_EXP(10),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_FPO_EXP(9),
      S01 => GRLFPC2_0_FPO_EXP(8),
      S10 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN21_LOCOV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un31_locov: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_FPO_EXP(10),
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPO_EXP(9),
      S11 => GRLFPC2_0_FPO_EXP(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN31_LOCOV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(3),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(43),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_0_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_1_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_1_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_2_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_2_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_2_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_3_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_3_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_3_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_3_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_4_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_4_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_4_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_4_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_5_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_5_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_5_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_5_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_6_2x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_6_3x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore_0: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore_1: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore_2: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore_3: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore_4: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_1,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un2_notdecodedunimp_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(64),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(66),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un3_notdecodedunimp: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un3_notdecodedunimp_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(67),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un3_notdecodedunimp_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un4_notresetorunimp: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(66),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN4_NOTRESETORUNIMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_status_1_6x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STATUS_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_un1_temp: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_un7_u_rdn_n: OR2A port map (
      A => GRLFPC2_0_R_FSR_RD(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN7_U_RDN_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_un20_u_rdn_0: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
      B => GRLFPC2_0_R_FSR_RD(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_8_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8_CM8I(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN7_U_RDN_N,
      S10 => GRLFPC2_0_FPI_LDOP_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_8_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(9),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8_CM8I(9),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_8_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_8_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_10_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_10(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_aregxorbreg: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un1_grfpus: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN1_GRFPUS);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un4_aregsign_sel: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un4_aregsign_sel_0: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un4_aregsign_sel_0_0: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un5_temp: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN5_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un10_aregsign_sel_m: XA1 port map (
      A => GRLFPC2_0_OP2(63),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(0),
      C => GRLFPC2_0_FPI_LDOP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN10_AREGSIGN_SEL_M);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_togglesig: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_FPI_LDOP_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_togglesig_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un1_u_snnotdb: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => GRLFPC2_0_FPI_LDOP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un2_sigtaf38_37: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN2_SIGTAF38_37);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un12_u_snnotdb_1: AND3C port map (
      A => GRLFPC2_0_FPI_LDOP_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      C => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un58_sctrl_new: AND4B port map (
      A => cpi_d_inst(12),
      B => cpi_d_inst(8),
      C => cpi_d_inst(11),
      D => cpi_d_inst(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN58_SCTRL_NEW);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp2_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(71),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN5_S_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp_1_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(73),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(73),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_1_CM8I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(72),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp_1_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(74),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_2(77),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_CM8I,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC,
      S11 => GRLFPC2_0_FPI_LDOP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_1_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_6: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_7: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_8: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_9: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_10: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_11: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_12: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_13: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_14: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_15: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_cm8i: CM8INV port map (
      A => GRLFPC2_0_FPI_LDOP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_temp: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(72),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(76),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un3_preventswap: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un5_notshiftcount1: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN5_NOTSHIFTCOUNT1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un17_srtosticky_0: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(11),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un17_srtosticky_1: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(9),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un17_wqstsets_n: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN5_NOTSHIFTCOUNT1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un42_conditional: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAINFNAN,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0(3),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(5),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4_N,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL_CM8I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un42_conditional_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_1: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_2: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_3: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_3_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_4: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1_5: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS_N,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_UN2_TEMP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_0: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS_N,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_UN2_TEMP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_1: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS_N,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1_CM8I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_UN2_TEMP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_1_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_1_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_un2_temp: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_UN2_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTBINFNAN_N,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_N,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_CM8I(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_6_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_5x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4(5),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_CM8I(5),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0_N(5),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_7x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN21_LOCOV,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN31_LOCOV,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_9x: OR3 port map (
      A => GRLFPC2_0_FPO_FRAC_0(54),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_0_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0_CM8I(3),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_0_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_0_n_5x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0_N(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4_5x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4_n_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4_N_CM8I(6),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4_N(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4_n_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4_N_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_6_6x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_6_CM8I(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4_N(6),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_6(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_6_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_6_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_conditional_6x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(9),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_a2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_A2_CM8I(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_253,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_275);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_a2_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_A2_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_a7_0_0_n_0x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_A7_0_N(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_a7_1_0x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_265);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_a7_2_0x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_266);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_o2_0_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_O2_0_CM8I(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_253);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_0_o2_0_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_0_O2_0_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_256,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_248,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_254,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_CM8I(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_243);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_0_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_265,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0_CM8I(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_0_3x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_0_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_1_2x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_245_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_2_3x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_245_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(3),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a2_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A2_CM8I(3),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_276);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a2_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A2_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a7_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_254,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_276,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_269);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a7_3x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_254,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_276,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_270);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a7_0_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_CM8I(2),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a7_0_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_1_CM8I(1),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a7_0_1_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_a7_0_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_A7_0_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_o2_1x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_248);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_o2_3x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_254);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_31_i_o2_0_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_256);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_0_sqmuxa_1_0: CM8 port map (
      D0 => GRLFPC2_0_FPI_LDOP_1,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3067,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_0_SQMUXA_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_3x: CM8 port map (
      D0 => GRLFPC2_0_OP2(51),
      D1 => GRLFPC2_0_OP2(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_26x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => rfo2_data2(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_27x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => rfo2_data2(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_28x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => rfo2_data2(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_29x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => rfo2_data2(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_30x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => rfo2_data2(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_31x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11),
      B => rfo2_data2(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_33x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_34x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_35x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_36x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_37x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_38x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_39x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_40x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11),
      B => rfo2_data2(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_41x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_42x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_43x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_44x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_45x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_46x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_49x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11),
      B => rfo2_data2(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_50x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data2(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_51x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data2(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_52x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data2(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_53x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data2(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_84x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data1(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_85x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data1(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_86x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data1(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(86));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_87x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11),
      B => rfo2_data1(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(87));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_88x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(88));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_89x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(89));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_90x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(90));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_91x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(91));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_92x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(92));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_93x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(93));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_94x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(94));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_98x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      B => rfo2_data1(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(98));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3713);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3714);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3715);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I(7),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3716);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3717);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I(9),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3718);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1_0_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_fprf_dout1_m_63x: AND2 port map (
      A => GRLFPC2_0_OP1(63),
      B => GRLFPC2_0_FPI_LDOP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPRF_DOUT1_M(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_4: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(244),
      fci => NN_4,
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(0),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_7: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(235),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(9),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(9),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_10: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(239),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(5),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(5),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_13: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(243),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(1),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_16: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(234),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(10),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(10),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_19: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(238),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(6),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(6),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_22: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(242),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(2),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(2),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_25: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(233),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(11),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(11),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_28: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(237),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(7),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(7),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_31: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(241),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(3),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(3),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_34: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(232),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(12),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(12),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_N_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_37: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(236),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(8),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(8),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_0_0_I_40: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(240),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(4),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(4),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_10,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_232);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_0: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_1: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_7: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_7_CM8I,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_7_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_7_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_9: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_248,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_9_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m1_10: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_0(3),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_7,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m5: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M5_CM8I,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M5_CM8I,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_10,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M1_9,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_270,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_31_I_2(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SLCONTROL(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m5_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_M5_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(5),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(5),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N(5),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1372,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_675,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(7),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(7),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N(7),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1344,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_20x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1262,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(21),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_30x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1194,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(30),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N(30),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_464,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4887_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1128,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_36x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(36),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(36),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N(36),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10(36),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1097,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(40),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1097,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_51x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10(51),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N(51),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(51),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_61x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(61),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(61),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N(61),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(4),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_N(4),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(4),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1025,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1450,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1477,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1097,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5057,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_24x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1643,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_914,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1641,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_27x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18(27),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_N(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(27),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(27),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_773,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_30x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1477,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1197,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_31x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19(31),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4455_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_1(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_32x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(32),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N(32),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(32),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(32),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_34x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4056,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1477,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1444,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_48x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(48),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_N(48),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_49x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_478_I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4977_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_992,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_53x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(53),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(53),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(53),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_54x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(54),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4885_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(54),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_55x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19(55),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N(55),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(55),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_57x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20(57),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21(58),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_N(58),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1324,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_4x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3989,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3988,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_18x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4610_1,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4181,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4303,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(27),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_29x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4410,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4396,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(29),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4410,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_1(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(58),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_0_0(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5285,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5285,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5285,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(59),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_62x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5406,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5406,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_0_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3926,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_4x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3985_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5193_I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_1_N(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_1(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_57x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_1_N(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_1(58),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(58),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(58),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5179,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_1_55x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4962_1,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5193_I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4959,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_1_tz_tz_55x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_20_0(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_TZ_TZ(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_1(0),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3937,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3938,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3990,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3990,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3990,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_9_1(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_CM8I(55),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4569_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_n_19x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_N_CM8I(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_N(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_n_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_15_0(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_N_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_2_tz_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4719,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_TZ(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_0(6),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4176_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4304,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_TZ_TZ(55),
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I(55),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4977_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5141_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_1_1(62),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5413,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I(62),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_1_1(62),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5407,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5402,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_cm8i_62x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_CM8I(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_n_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_N_CM8I(29),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0(29),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4402,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(29),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4409,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_N(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_n_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4412,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_N_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_tz_n_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_TZ_N_CM8I(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4649_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_TZ_N(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_3_tz_n_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_1_0_N(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_TZ_N_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4182_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I(18),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_1_N(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_13_1(32),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I(32),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4525_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I(58),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_11_0_N(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4528_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_n_0x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(0),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3935,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_n_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N_CM8I(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_n_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N_CM8I(28),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N_CM8I(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4375_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4374,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4371,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_n_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_4_n_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4377,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3936,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4043,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4182_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I(18),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4370,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_1_0(28),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4373,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5218,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_0_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4462,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_4_1(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_5_n_62x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5403,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_N(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_4x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3969,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4026,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4056,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4046,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4470_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_7_0(59),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(59),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I(59),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5393,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(62),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5405_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_5_1(62),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I(62),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_0_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4471,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4458,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_cm8i_62x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_0_0(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_CM8I(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_n_32x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_N_CM8I(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4545_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4541,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_N(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_6_n_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_N_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3969,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4679,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4685,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_55x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_CM8I(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4966_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4981,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5290,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_22_1(59),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5272,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_n_6x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N_CM8I(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_n_32x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N_CM8I(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_0(32),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4531,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4540,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_n_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4055_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_7_n_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4502,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4465,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4430,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4502,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4465,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_32x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4533,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4543,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4535,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4677,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_52x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(52),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4756_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4765,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4763,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_53x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4765,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_0(53),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(54),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_19_0(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4127_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_1_N(54),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_59x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5271,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_4_0(59),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4962_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_21_0(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4708,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_1(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4890_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_10_1(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I(4),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3983,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3987,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3990,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_6x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5410,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4052,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4321,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_27x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1349,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_6546,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4314,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_58x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I(58),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(58),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5132_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3981,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_n_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_tz_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_TZ_CM8I(18),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_TZ(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_8_tz_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_TZ_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_6x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4061,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_18x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1(18),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4545_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_11_1(19),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4225,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_19_0(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4225,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4306,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4292,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_32x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(32),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4564,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4536,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1262,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4184_1,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4683,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_11_1(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4683,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_52x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4753,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4761,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4749,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_54x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4887_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4962_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_1(59),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(59),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_0_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4502,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_0_CM8I(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_0_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_2_1(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_0_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4710,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_0(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4513_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_n_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N_CM8I(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N_CM8I(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_n_53x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4766_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4802,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4829,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4832,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_9_n_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_0(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3991,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4055_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4171,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4179,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_13_0(19),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4239,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_5_0(19),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4239,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1117,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_0_0(32),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4522,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_17_1(48),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4678_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_0(48),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_52x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_0(52),
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4748_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I(52),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4824,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4811,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4830,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_1(54),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_TZ_N(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_0(57),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(57),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5107,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4750,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_10_n_4x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1257,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10_N(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4(18),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4184_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_TZ(18),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(18),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_23_1(31),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4460,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1197,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_48x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4691,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4686,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4680,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4784,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_0(52),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_CM8I(52),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4784,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4759,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4755,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_53x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_CM8I(53),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4831,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4817,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4886,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_0(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5134,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_19_0(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5133,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4766_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4802,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_n_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_N_CM8I(27),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4289,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_1(27),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4710,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_10_0(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_N(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_11_n_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11_N_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_4x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3984,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I(4),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(4),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3992,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3979,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_27x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4311,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4319,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4316,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_6545,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_31x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_0(31),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4675,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4687_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_TZ(48),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4681,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4674,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4760,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_14_0(52),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4757,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4769,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_53x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4825,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4823_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4828,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4820,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_54x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4893,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4889_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4904,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4758,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_55x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4979,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4979,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4979,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4835,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4899,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_n_57x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_17_1(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5136,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_n_59x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_20_0_N(59),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N_CM8I(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_12_n_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5284_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_19x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_0(19),
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(27),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_1(27),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4324,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(31),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13_CM8I(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_1(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4896,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(57),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5097_I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5132_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5131,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5124,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_59x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5292,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5282,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5270,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_13_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4226,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_1(19),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4224,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_31x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3945,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4428_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4961,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4972,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4960,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_1_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_0(31),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4449,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_1_0(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4467,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4480,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_n_48x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(48),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_N(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_14_n_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4678_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5182,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5201,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14_N(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_19x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4245,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4247,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4246,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4235,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_32x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4530,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I(32),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6_N(32),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4537,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_0(57),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I(57),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5137,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5222_1,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(58),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5208_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4538,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5169,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_15_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5205,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_16_6x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4058,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4045,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_16_53x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(53),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(53),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4822,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4819,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_16_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4955,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_18_1(55),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_1(55),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_16_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5122,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_15_0(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5182,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5127,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5139,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_16_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5214,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16_CM8I(58),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5212,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_16_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5207,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_19x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4228,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_CM8I(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2_N(19),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4242,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4237,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_52x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(52),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4747,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4751,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4758,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_54x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(54),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(54),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_2(55),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_12_0(55),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4975,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4963,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_59x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5289,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_CM8I(59),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5279_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5287,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5276,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5273,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_n_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_N_CM8I(58),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5223_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5206,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5204,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_N(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_17_n_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5215,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_N_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_18_27x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4302,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_CM8I(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(27),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(27),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_18_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_1(55),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(55),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_CM8I(55),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_18_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4321,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_18_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_18_n_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8_N(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_N_CM8I(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7_N(6),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1151,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_N(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_18_n_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4041,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_N_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_6x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(6),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4040,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4053,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_31x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(31),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_N(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_CM8I(31),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9_0(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_55x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(55),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4978_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_CM8I(55),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4964,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4969,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4967,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_n_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_N_CM8I(52),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(52),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4752,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_N(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_19_n_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(52),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_N_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_20_52x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(52),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(52),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_989,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_20_57x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(57),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(57),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_20_n_19x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(19),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(19),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_20_n_55x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(55),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_922,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_20_n_59x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17(59),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(59),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_21_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(19),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4227_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I(19),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(19),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_21_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I(58),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_17_N(58),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_21_59x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_14(59),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I(59),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12_N(59),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(59),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_21_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4210,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_21_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_21_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3945);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_28x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_4x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_18x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_53x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_62x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5413);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_0_18x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_0_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_0_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_0_0_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_27x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_28x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4382);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_29x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4417);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_0_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_0_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_1_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_1_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_1_1_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_2_18x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4545_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_2_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_2_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_2_58x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_2_0_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_3_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_3_0_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_4_28x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_4_29x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4421);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_5_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_5_52x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4784);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_5_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5284_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_5_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5302);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_5_62x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5418);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3923_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_19x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4260);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_0_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_0_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_1_0x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_1_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_6_1_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_7_19x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_7_27x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_7_29x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_7_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4708);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_7_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_7_0_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_54x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5164);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_0_54x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_0_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_0_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_8_1_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_9_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4710);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_9_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5165);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_9_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_9_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_9_0_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_9_0_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_31x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_32x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_52x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_53x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_58x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5246);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_0_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_1_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_1_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_10_2_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_27x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4347);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_32x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5410);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_0_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_1_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_11_2_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_12_32x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4564);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_12_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_12_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_12_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_13_6x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4081);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_13_27x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_13_31x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4502);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_13_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5169);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_13_58x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_13_0_58x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_14_19x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4269);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_14_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5004);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_16_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_16_0_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_16_1_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_16_2_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_18_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4719);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_19_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_19_0_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a2_20_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4699);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a7_0_29x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a7_0_2_29x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4408_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a7_1_29x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4417,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4409);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a7_2_29x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4398,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4410);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a7_4_29x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4412);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_CM8I(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3935);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_28x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_CM8I(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4370);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_0_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3936);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_0_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4382,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_CM8I(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4371);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_0_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_0_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_1_0x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3931,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3937);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_1_0_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_1_0(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_2_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_2_CM8I(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3938);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_2_28x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_2_CM8I(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4382,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4373);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_2_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_2_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_2_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_2_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_3_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_CM8I(28),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4374);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_3_0_0x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_3_1_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_3_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_4_1_28x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4375_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_5_28x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_5_0_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_5_1_0x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_5_2_28x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_6_28x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4377);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a9_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_62x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5390,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4129_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_CM8I(62),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4129_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_0_0_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_0_0(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_1_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_1_1_62x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_1_1(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_2_62x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4428_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5402);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_3_62x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5403);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_5_1_62x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5405_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_5_1_0_62x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_5_1(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_6_62x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5418,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5406);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_7_62x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5418,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5407);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a10_cm8i_62x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A10_CM8I(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_1_18x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4171);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_1_2_18x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_4_1_n_18x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_1_N(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_5_18x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_6_1_18x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4176_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_9_18x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4176_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4179);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_11_18x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4181);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_12_1_18x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4182_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a17_14_1_18x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4184_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_4x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_0(4),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3979);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_0_0_4x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_1_4x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3968,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3981);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_2_1_n_4x: OR3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_1_N(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_3_4x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_2,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3983);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_3_1_4x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_4_4x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3965_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3984);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_5_1_4x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3985_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_6_1_4x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_7_4x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3987);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_8_4x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4018,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3988);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_9_4x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4018,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3989);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_10_4x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3990);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_11_4x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3991);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_12_4x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_12_0(4),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3992);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a18_12_0_4x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_12_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_0_0_0_32x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_0_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_1_32x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_CM8I(32),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4530);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_1_0_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4528_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_1_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_2_32x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4520,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4531);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_3_0_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_4_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_4_CM8I(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4533);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_4_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_4_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_5_32x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4513_I,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_5_1_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_6_32x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4535);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_7_32x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4977_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4536);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_8_32x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3923_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4537);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_9_32x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3923_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4538);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_11_32x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4540);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_12_32x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5222_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4541);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_12_1_32x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5222_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_13_1_32x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_13_1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a20_14_32x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4543);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_48x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4710,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_0_48x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673_1,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_CM8I(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_0_53x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4810,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4817);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_0_1_53x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_0_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_1_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4111_1,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_CM8I(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4674);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_1_0_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4672_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_1_0_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_0_CM8I(53),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_0(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_1_0_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_0_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_1_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_2_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_CM8I(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4675);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_2_53x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_CM8I(53),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4819);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_2_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_2_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4699,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_3_53x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_CM8I(53),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4820);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_3_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_4_48x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4677);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_5_53x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4822);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_5_0_48x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_5_1_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4678_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_6_48x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4719,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4708,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_6_CM8I(48),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4719,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4679);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_6_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_6_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_6_n_53x: OR4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5193_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4823_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_7_48x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4699,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4680);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_7_53x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4824);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_8_48x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_CM8I(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4708,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4681);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_8_53x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4408_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4825);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_8_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_9_0_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4649_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_9_1_53x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_1(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_10_48x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4708,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4683);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_10_1_53x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_11_53x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4828);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_11_1_48x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_11_1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_12_48x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4685);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_12_53x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4829);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_13_48x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4686);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_13_53x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4830);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_14_53x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4831);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_14_1_48x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4687_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_15_53x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4832);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_16_1_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_16_1_0_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_17_1_48x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_17_1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_18_48x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4691);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a21_18_53x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4835);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4018,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4081,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_CM8I(6),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4081,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4040);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_0_6x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4032,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4041);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_0_54x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4886);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_1_1_54x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4887_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_2_6x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_CM8I(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4043);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_2_54x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888_1,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_CM8I(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_2_1_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_2_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_2_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_3_n_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_N_CM8I(54),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4889_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_3_n_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_N_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_4_6x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4045);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_4_n_54x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5179,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4890_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_5_6x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4046);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_5_1_54x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_6_0_54x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4892_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_0(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_6_1_54x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4892_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_7_54x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_CM8I(54),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_1_0_N(54),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4893);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_7_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_9_1_n_54x: OR3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_1_N(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_10_54x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4896);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_11_6x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4052);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_11_1_54x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_12_6x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4081,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4053);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_13_54x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4899);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_13_0_6x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_14_1_6x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4055_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_14_1_54x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5179,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_15_6x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4056);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_15_54x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_16_1_54x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_17_6x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4058);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_17_54x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4903);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_18_54x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4904);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_19_0_54x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_19_0(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_19_1_54x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4127_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_20_6x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4061);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_20_1_0_n_54x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_1_0_N(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_n_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_N_CM8I(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4885_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a23_n_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5284_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_N_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4347,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4285,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_CM8I(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4302);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_52x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4744,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5302,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4747);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_0_27x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4303);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_0_n_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4748_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_1_27x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4802,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4304);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_1_52x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4739,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4749);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_2_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_2_CM8I(52),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4750);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_2_1_27x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_2_2_27x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_2_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_2_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_3_27x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_3_CM8I(27),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3923_I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4306);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_3_52x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4616_1,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4751);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_3_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_3_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_4_52x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1003,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4752);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_4_1_27x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_5_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_5_CM8I(52),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4753);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_5_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_5_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_6_0_52x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_6_1_27x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4699,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_7_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_7_CM8I(27),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_6545);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_7_52x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4428_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4755);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_7_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_7_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_8_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_8_CM8I(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4311);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_8_1_52x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4756_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_8_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_8_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_9_27x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_6546);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_9_52x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4757);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_10_52x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4758);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_10_0_27x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_10_0(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_11_27x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4314);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_11_52x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4759);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_12_52x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4760);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_13_27x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4316);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_13_52x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4761);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_14_0_52x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_14_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_15_52x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5302,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4763);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_16_27x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4319);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_17_27x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5164,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_17_52x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4765);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_17_1_27x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_18_27x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4710,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4321);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_18_1_52x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4766_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_19_0_52x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_21_27x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4320_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4324);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_21_52x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4616_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4769);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a24_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4224);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_59x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_CM8I(59),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4839,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5270);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_0_19x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_0_CM8I(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4225);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_0_59x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5302,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5271);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_0_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_0_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_1_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_1_CM8I(19),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4269,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4226);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_1_59x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5272);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_1_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_1_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_2_59x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5273);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_3_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_3_CM8I(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4228);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_3_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_3_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_4_19x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_4_0_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_4_0(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_4_1_19x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_5_59x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5276);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_5_0_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4260,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_5_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_6_0_19x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_6_1_19x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4231_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_6_1_59x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_1(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_7_19x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_7_0_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_7_0(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_7_2_19x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4232_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_8_n_59x: OR4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5279_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_9_1_19x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4269,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_10_19x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4235);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_10_1_59x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_10_1(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_11_59x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5282);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_11_1_19x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_11_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_12_19x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4227_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4237);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_12_1_19x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4227_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4237_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_12_1_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5283_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_13_0_19x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4229_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_13_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_14_19x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4239);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_14_59x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5285);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_15_59x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_15_0_19x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3997,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_15_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_15_1_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_16_59x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5287);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_17_19x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4242);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_18_59x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5289);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_19_59x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5164,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5290);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_19_0_19x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4260,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_19_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_20_19x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4245);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_20_0_n_59x: OR3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_20_0_N(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_21_19x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4246);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_21_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_21_CM8I(59),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5292);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_21_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_21_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_22_19x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4247);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_22_1_59x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_22_1(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a25_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_57x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5122);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_58x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4231_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_CM8I(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5201);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_0_0_58x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_0_0(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_0_1_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_1_57x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5110,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5124);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_1_58x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5193_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_1_1_58x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_2_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5246,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_CM8I(58),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5204);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_2_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_2_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_3_58x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5205);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_3_0_57x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_4_57x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5169,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5127);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_4_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5206);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_5_58x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5246,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5207);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_5_1_n_57x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_1_N_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_1_N(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_5_1_n_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_1_N_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_6_1_57x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5101_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_6_n_58x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_N_CM8I(58),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5208_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_6_n_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_N_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_7_57x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5164,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_7_1_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_1(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_7_2_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5130_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_8_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_8_CM8I(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5131);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_8_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5164,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_8_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_9_58x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_9_1_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5132_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_10_57x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_10_58x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5179,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5212);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_11_57x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5134);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_11_0_n_58x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5412,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_11_0_N(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_12_58x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5214);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_12_1_57x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_13_57x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5136);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_13_58x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5211_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5215);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_14_57x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5091,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5137);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_15_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5165,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_15_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_15_1_58x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5229,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5217_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_16_57x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5182,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5139);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_16_58x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4305_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5218);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_17_1_57x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5301,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_17_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_18_2_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5141_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_19_0_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4528_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_19_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_20_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_20_1_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_21_1_58x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5223_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_22_58x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_22_1_58x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5224_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a26_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_55x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5004,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4955);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_0_1_55x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_0_n_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_N_CM8I(31),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5405_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4455_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_0_n_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_N_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_1_0_31x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4470_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_1_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_1_0_55x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_1_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_2_1_31x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_2_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_2_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_2_1_0_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_3_31x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4443,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_3_0(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4458);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_3_55x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4939_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5419_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4959);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_3_0_31x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_3_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_4_55x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4938,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4960);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_4_1_31x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_4_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_5_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_0,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4460);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_5_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231_1,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_5_CM8I(55),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4961);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_5_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_5_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_6_0_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_0_CM8I(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4260,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_6_0_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_0_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_6_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4962_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_7_31x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_478_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4462);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_7_55x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4963);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_8_55x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4964);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_9_1_55x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_9_1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_10_31x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_10_CM8I(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4465);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_10_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4966_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_10_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_10_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_11_55x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4967);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_12_31x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4428_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4467);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_12_0_55x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_12_0(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_13_55x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4969);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_14_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_14_1_0_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_15_1_31x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4470_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_16_31x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4471);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_16_55x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4972);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_17_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_18_1_55x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_18_1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_19_55x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5004,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4975);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_20_0_55x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_20_0(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_21_0_31x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_21_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_21_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4977_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_22_n_55x: OR4D port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4978_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_23_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4979);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_23_1_31x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_23_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_23_1_55x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_25_31x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5233,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4480);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_a28_25_55x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4981);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_12(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_8(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4756_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_7(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1607,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_16(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_13(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_15(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4018);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(19),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4210);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4285);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4395);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4520);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4739);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(57),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5107);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_0_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4443);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m2_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_m28_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5399_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4938);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_1x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_2x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1304,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(8),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(14),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_33x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_627,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(42),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(43),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_989,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4618_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_n_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_53x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_0_48x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_0_53x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_0_62x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5410,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5390);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_0_0_48x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_1_53x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o2_2_53x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o7_29x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4424,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4396);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o7_0_29x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4395,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4398);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o7_2_29x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4421,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4402);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o9_1_0x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3945,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3926);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o9_3_0x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4124_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3931);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o10_62x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o10_0_62x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o10_0_0_62x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o10_0_1_62x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o10_3_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5393);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o17_2_18x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o17_2_0_18x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o18_0_4x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o18_0_0_4x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o18_3_4x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3968);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o18_4_4x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3969);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o20_0_32x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o20_0_0_32x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o20_4_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4564,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4522);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o20_5_n_32x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4563,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4525_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o21_3_53x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o21_3_0_53x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o21_3_1_53x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o21_4_53x: OR2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4802);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o21_7_53x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_478_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4810);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o21_8_53x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4811);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_0_54x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_0_0_54x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_0_1_54x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_3_6x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_3_0_6x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_5_6x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4026);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_6_6x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4032);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_8_54x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o23_8_0_54x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o24_1_52x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o24_2_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5422,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4289);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o24_4_27x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4292);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o24_6_52x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4744);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_0_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_2_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_2_0_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_3_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_3_0_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_3_1_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_3_2_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o25_5_59x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5256);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_0_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_0_58x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_0_0_58x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_1_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_1_58x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_1_0_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_1_1_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_1_2_57x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_2_58x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5179);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_3_57x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5167,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5165,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5091);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_3_58x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_3_0_58x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_3_1_58x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_4_58x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5182);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_5_57x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_5_0_57x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_5_1_57x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_11_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_11_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5110);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o26_11_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_11_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O28_CM8I(31),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4430);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_0_55x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_0_0_55x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_1_55x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_1_0_55x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_1_1_55x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_1_2_55x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_3_31x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4449);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_o28_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O28_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_4x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3965_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_6x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_32x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4513_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_48x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_53x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_54x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_55x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4939_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_57x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_58x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_62x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_0_48x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4649_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_0_52x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4428_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_0_54x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_0_57x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_0_58x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5193_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_0_62x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_1_53x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_478_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_1_55x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4569_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_1_57x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5101_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_2_27x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_2_57x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5097_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_2_0_27x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_0_x2_3_27x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3923_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0(7),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(7),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_12x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1605,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1304,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_26x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1077,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4673_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(34),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN5_S_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_36x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1600,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1502_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1092,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(41),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1092,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_1(7),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(50),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_0_5x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1639,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_0_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1539,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0_CM8I(7),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_0_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_1_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1480,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1517,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_2_n_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_2_N_CM8I(17),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_2_n_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_2_N_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_440_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_n_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N_CM8I(3),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1391,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_n_30x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1195,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_1_n_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1493,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_5x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1302,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1300,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_23x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1256,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1257,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1247,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I(25),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_26x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4888_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_30x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1480,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_34x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(34),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1133,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_36x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1116,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_38x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1103_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I(38),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_49x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1523,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1523,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1664,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1108,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_cm8i_61x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_CM8I(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_10x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1486,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1485,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_15x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1641,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1302,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_37x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1110_N,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1109_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I(37),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1107,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1418,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I(39),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1101,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_464,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I(41),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1111,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1100,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_2_n_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_15x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_761,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1276,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1300,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1643,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1151,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1113,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1448,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I(36),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1113,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1486,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I(37),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1104,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I(38),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1104,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_49x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_TZ(49),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_50x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1477,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_61x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_765,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1103_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_n_17x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1298_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1566,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_N(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_3_n_25x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1245,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1391,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_N(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_5x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I(5),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1244,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I(25),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1244,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_34x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1014,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1010,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1582,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_n_44x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_500,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_N(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_4_tz_49x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1637,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_TZ(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_989,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_989,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_CM8I(7),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1151,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1346,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1666,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1084,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(49),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_61x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1666,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_0_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_n_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N_CM8I(12),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1324,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1256,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_n_13x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1317,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_n_33x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N_CM8I(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_n_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_5_n_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1656,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_12x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_1(17),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_482,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_34x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_CM8I(34),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_38x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(38),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1101,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1100,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_440_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_n_3x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N_CM8I(3),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1389_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1276,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_n_7x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1093,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1352,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1543,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_n_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N_CM8I(26),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_611,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1027,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_n_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1650,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_6_n_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_482,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_7x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1637,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1300,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_690,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(26),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_49x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(49),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1656,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4598_1,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1656,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5289,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1003,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_0_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(7),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1493,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1349,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1092,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_n_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N_CM8I(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N_CM8I(17),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_n_33x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1609,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_n_61x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(61),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_7_n_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1324,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I(5),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_1(7),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_500,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(13),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1605,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4237_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1310,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(33),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_914,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_34x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1132,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(34),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1135,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1117,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_663,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4973_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I(36),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1117,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(51),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(61),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I(61),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_3_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1647,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_8_cm8i_61x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1493,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8_CM8I(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1312,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1315,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_25x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303_0,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3991,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_589,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(33),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(34),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_CM8I(34),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_36x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_589,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(51),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4756_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(61),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1582,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_768,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_n_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N_CM8I(5),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(5),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1371,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_n_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N_CM8I(50),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_501,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(50),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_n_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_0(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_9_n_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1084,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_CM8I(36),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1607,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(36),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(50),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_614,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_621,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_51x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_n_13x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N(13),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1448,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_0(13),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N_CM8I(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_n_17x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N_CM8I(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_N(17),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_507,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_n_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1607,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_10_n_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1276,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_13x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1045_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_17x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1_1(17),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_CM8I(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_N(17),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_482,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_590,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1148,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1141,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1298_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_CM8I(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(49),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(49),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1656,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_11_n_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4(25),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_690,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_N(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_12_25x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(25),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12_CM8I(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3_N(25),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(25),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1243,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_12_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_614,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1664,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_997,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_993,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_12_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_12_n_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6(34),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12_N(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_13_13x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1311_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1609,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_13_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(34),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4380,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(34),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_13_49x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(49),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13_CM8I(49),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1018_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1025,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_621,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_13_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1027,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_14_n_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N_CM8I(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N_CM8I(49),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(49),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_14_n_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1029,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_15_n_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N_CM8I(36),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(36),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_15_n_51x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N_CM8I(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1609,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_0(51),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_15_n_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_15_n_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_15_N_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_16_n_33x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7_N(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_16_N_CM8I(33),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N(33),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(33),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_16_N(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_16_n_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_16_N_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_17_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(33),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_17(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_17_n_13x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_675,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_8(13),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_17_N(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_18_13x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13(13),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_18_CM8I(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N(13),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1306,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_18(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_18_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_18_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_7x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1543);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_16x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5299,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1485);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_33x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1609);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_37x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1414,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1637,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1418);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_49x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1445,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1607);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_53x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_58x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_3x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1650);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_CM8I(16),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_0(62),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_663,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1486);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_17x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1517);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_24x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1592);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_39x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_42x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1539);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_53x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_0_n_3x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_N(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_1_42x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_1_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_0_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_27x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1601);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_33x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1445);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_50x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_51x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_53x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1477);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_58x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1414);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_61x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_0_58x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1526_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_1_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_17x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1566);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_24x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1572);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_33x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1643);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_51x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1656);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_0_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_2_0_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1600);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_51x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1664);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1500);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_56x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1450);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_57x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_3_0_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_0(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_17x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1588);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_31x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1639);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_55x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1471);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1605);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_4_58x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1448);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_5_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_5_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_5_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4385,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_5_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_5_0_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_5_1_17x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1502_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_6_31x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_6_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_6_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_6_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_6_62x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_7_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_7_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_8_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_8_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_8_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1493);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_8_0_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_9_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_9_59x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1444);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_9_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_9_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_10_59x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_10_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1455);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_11_59x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_11_61x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1523);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_12_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_13_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1647);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_13_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_13_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_13_62x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5249,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_14_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_14_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1480);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_14_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1582);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_14_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_15_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_15_61x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1641);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_16_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1666);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a2_28_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1637);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1445,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1371);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_667_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1346);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_13x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1435,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1306);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_20x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1450,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1262);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_23x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1256);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_25x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1243);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_33x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1141);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_39x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1100);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_40x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1097);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_41x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1092);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_46x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1077);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1641,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_765);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_5x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1419,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1372);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_9x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1344);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_14x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1304);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_15x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1302);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_17x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4158,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4792_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_23x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1257);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_25x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4032,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1244);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_30x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1194);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_36x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4408_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1113);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_38x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1104);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_39x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1647,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1101);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_41x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1093);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_45x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_50x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1010);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_51x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_992);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_0_13x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_1_17x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1296_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_2_17x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1601,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_0_n_37x: OR2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1110_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_3x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1445,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1391);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_12x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1525,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1324);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_25x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5016_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1245);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_30x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5203_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1195);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_37x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1111);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_44x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_51x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5054,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_993);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_61x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_0_13x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_0_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_1_44x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1082_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_1_1_61x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5177,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_7x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1349);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_28x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1211);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_34x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1132);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_35x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1128);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_61x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_768);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_0_25x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_0_50x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_2_1_17x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1298_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_13x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4648_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1310);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_25x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4023_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1247);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_30x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1197);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_34x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1639,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1116);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_38x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1107);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_44x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1084);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_3_0_5x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_3_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_4_17x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1450,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1300);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_4_36x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1117);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_4_38x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1523,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1501,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1108);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_4_44x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1480,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_4_50x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4887_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1014);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_4_1_13x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1311_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_7x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1352);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_13x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1312);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_34x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1135);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_51x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_5_0(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_997);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_61x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_0_51x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5168,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_5_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_5_1_61x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_771_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_6_33x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4957_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1148);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_6_49x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1025);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_6_51x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7_13x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0(13),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1314);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7_59x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4507,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7_61x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1452,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1524,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_773);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7_62x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_761);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7_0_13x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_7_0_49x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_8_13x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1315);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_8_49x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1027);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_8_51x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1474,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_8_53x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1475,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_954);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_9_33x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1458,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1600,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1151);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_10_13x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1479,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4789,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1317);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_10_49x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1420,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1029);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_11_19x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1276);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_11_48x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4970_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_11_51x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5253,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1003);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_11_1_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_12_1_48x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1045_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_15_55x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4897_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_914);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_22_52x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1647,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_989);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_23_55x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1491,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4958_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_922);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_n_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4598_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1389_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_n_37x: OR3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4437_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1109_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_n_38x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_N_CM8I(38),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1103_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_n_49x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_N_CM8I(49),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1448,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1444,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1018_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_n_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_N_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_a12_n_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_N_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1635,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1428,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(51),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_cm8i_61x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_773,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_CM8I(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_0_47x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4612,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4603,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_0_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4843,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5286_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_0_tz_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_TZ_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_TZ(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_0_tz_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_TZ_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_1_n_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_1_N_CM8I(47),
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_1_N(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_1_n_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_1_N_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_2_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_1_0(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4099,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4871,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_2_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2_CM8I(60),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5093,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_2_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_4_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4125_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4113,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4_CM8I(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_4_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4618_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4616_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5087,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_4_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5040,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_4_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5344,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5344,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5344,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_4_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_5_11x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_5_CM8I(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_5(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_5_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_5_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_6_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_23_0(56),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_CM8I(56),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_6_60x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_10_0(60),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_CM8I(60),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_6_0_60x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_3_0(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5326,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5357,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5342,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_0(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_6_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_6_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_8_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_8_CM8I(47),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1637,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_8(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_8_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_8_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_9_11x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_3_0(11),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_9_CM8I(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4534_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4123,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4133,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_9(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_9_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_9_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_10_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4122,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4227_1,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4122,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_10_CM8I(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_10(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_10_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5252,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_10_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_11_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4111_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_0(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_11_CM8I(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_11(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_11_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4124_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_11_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_12_56x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_CM8I(56),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5054,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5348_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_12_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(60),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_12_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_12_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_12_n_47x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4928,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_N_CM8I(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_2_0(47),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4594,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4601,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_N(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_12_n_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4966_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_N_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_13_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_8_0(11),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4118,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_5(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_13_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4609,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_TZ(60),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5346,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_13_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_19_0(11),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(11),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_9_0(11),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_47x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I(47),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_56x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5030,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(56),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6_0(60),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5348_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5353,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4099,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_14_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_15_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4127_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4129_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_15_56x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5042,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5038,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_15_n_60x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15_N_CM8I(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5350_N,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5339_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5337,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15_N(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_15_n_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5343,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15_N_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_16_11x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4117,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16_CM8I(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4115_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4126,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4134,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_16_47x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4620,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16_CM8I(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4599_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4615,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_16_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_10_1(56),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5039,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_16_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4116,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_16_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4605,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_17_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_4(47),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4598_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_0(47),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4610,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4602,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_17_56x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17_CM8I(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5055_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5045,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_17_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5048,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_18_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_11(11),
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4129_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_2(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_18_47x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18_CM8I(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12_N(47),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_18_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5051_1,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18_CM8I(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5057,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5062,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_18_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4606,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_18_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_19_47x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_8(47),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_CM8I(47),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_1_N(47),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(47),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4609,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_19_56x: OR4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12(56),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5036,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5046,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5044,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_19_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4596,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_19_n_60x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15_N(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_N_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5336_N,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5338,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_N(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_19_n_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_6(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_N_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_20_n_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_20_N_CM8I(60),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1093,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13(60),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_20_N(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_20_n_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_12(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_20_N_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_21_n_11x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18(11),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_9(11),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_21_N(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_22_n_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N_CM8I(11),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16(11),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_22_n_47x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4595,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_22_n_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_13(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_23_n_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N_CM8I(47),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17(47),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1211,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_23_n_56x: AND3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19(56),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_14(56),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_15(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_23_n_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_24_n_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_24_N_CM8I(56),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_4_0(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5024,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_17(56),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_18(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_24_N(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_24_n_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_16(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_24_N_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_47x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_0_47x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_0_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_0_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_0_0_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_1_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_2_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_0_3_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_1_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_1_0_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_1_1_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_2_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_2_0_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_3_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4227_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_4_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_5_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_5_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_5_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_5_0_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_5_1_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_6_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_6_0_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_8_60x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_8_0_60x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_9_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_9_0_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_9_1_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_11_47x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_12_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_12_0_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_12_1_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a2_12_1_0_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_0_60x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5337);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_0_0_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_0_CM8I(11),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_0_0_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_0_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_0_1_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4111_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_0_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_0_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_1_60x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1647,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5089,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5374,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5338);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_1_0_11x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5295,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_1_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_2_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5165,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_2_CM8I(11),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4113);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_2_1_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_2_1(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_2_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_2_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_2_n_60x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_2_1(60),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5339_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_3_0_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_3_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_3_0_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_3_0(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_4_60x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5380,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5341);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_4_n_11x: OR4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4115_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_5_11x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4116);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_5_60x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5321_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5342);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_6_11x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4093_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4117);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_6_60x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_667_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5343);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_7_11x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5418,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5244,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4118);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_7_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_7_CM8I(60),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5344);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_7_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_7_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_8_0_11x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4555,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_8_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_8_1_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_9_60x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5346);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_9_0_11x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_9_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_10_0_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_10_0(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_10_1_11x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4901_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_11_11x: AND4A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717_2,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4122);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_11_2_60x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5418,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5348_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_12_11x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4123);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_13_1_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4273_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4124_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_13_n_60x: OR4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5350_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_14_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_14_1_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_14_2_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4125_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_15_11x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4499,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4126);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_15_1_60x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5352_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_16_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5351_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5353);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_18_1_11x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4129_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_19_0_11x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_19_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_19_1_60x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_20_60x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5357);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_22_11x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4017,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5155,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_23_11x: AND4 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5163,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5161,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4134);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_n_60x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_N_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5336_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a26_n_cm8i_60x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5362,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_N_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_47x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4592,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4921,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4594);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_56x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3985_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_CM8I(56),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5036);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_0_47x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1045_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_0_CM8I(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4595);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_0_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_0_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_1_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5379,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_1_CM8I(47),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4596);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_1_56x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5038);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_1_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_1_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_2_56x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_2_CM8I(56),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5028,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5039);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_2_0_47x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4795,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_2_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_2_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4727,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_2_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_3_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_CM8I(56),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5040);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_3_0_47x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_0_CM8I(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_3_0_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_0_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_3_1_47x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4598_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_3_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_3_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_4_0_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4996,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_4_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_4_n_47x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4330,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5141_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4892_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4599_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_5_56x: XA1 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4887_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5042);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_6_47x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5234,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4986,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4601);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_6_56x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5071,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_6_1_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5043_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_7_47x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4697,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4602);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_7_56x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5387,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5016_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5044);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_8_47x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5178,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4603);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_8_56x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5045);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_9_56x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4562,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5046);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_10_47x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4569_I,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4605);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_10_1_56x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_10_1(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_11_47x: AND4C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4569_I,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4606);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_11_56x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5048);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_14_47x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4631,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4717,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4609);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_14_1_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5051_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_15_47x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4610);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_15_1_47x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4632,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4610_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_17_47x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4623,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4612);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_17_56x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1591_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5054);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_17_1_56x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1591_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_18_n_56x: OR3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5075,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5055_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_20_47x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4799,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5076,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4615);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_20_56x: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5057);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_21_1_47x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5388,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4616_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_23_0_56x: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4910,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_23_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_23_1_47x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4645,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4927,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4618_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_24_56x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5180,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_24_1_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5061_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_25_47x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4858,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4892_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4620);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_25_56x: AND4B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3959,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5001,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5231,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5062);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_a28_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_0_56x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_0_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5310_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_0_0_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_0_0_0_56x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_0_1_56x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_0_2_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5008_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_1_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_1_0_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o2_1_1_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_0_60x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5311);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_0_0_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_1_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_1_0_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_1_1_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_4_60x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5312,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5326);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o26_5_11x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5152,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4099);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_0_47x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_0_0_47x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4575_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_1_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5015);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_2_56x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_O28_2_CM8I(56),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5361,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5242,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5421,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5024);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_2_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_O28_2_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_4_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5082,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5028);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_6_56x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5013,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5030);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_o28_8_47x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4638,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4592);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_x2_56x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4094_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_x2_60x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_433_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_x2_0_56x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5016_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_x2_0_60x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_667_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_x2_1_60x: XNOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4581_I,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5321_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_i_x2_2_60x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4360_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_m2_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_M2_CM8I(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_627);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_m2_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_M2_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_34x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1497,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_36x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_663);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_52x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_0_32x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_611);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_0_50x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1417,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_501);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_0_52x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_0_56x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4262,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_1_47x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_1_52x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_1_58x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_1_0_58x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o2_4_60x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_488);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1482,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_N(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_5x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5143_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1468,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_482);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1276,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1650,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1300,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_678);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_922,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1441,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1077,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1601,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_507);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_24x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1500,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0(26),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(26),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_690);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_34x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1317,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4412,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1315,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(36),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1418,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0(39),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1471,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1107,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_464);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1085,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1476,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4061,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1444,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_500);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_50x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1471,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_507,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_621);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_51x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1440,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1449,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4698,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_614);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1433,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_761,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1425,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_CM8I(13),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_761,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_675);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_24x: OR3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1572,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0(24),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1592,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_646);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1431,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4372_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_449_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_CM8I(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4827_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4625,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_412,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1211,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5000,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3952_1,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_38x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3954,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1430,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5345_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_39x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1103_N,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1486,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_559);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_0_0_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5068,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1493,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5356_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0_0_CM8I(24),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5309,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_0_0_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5294,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0_0_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4689_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_0_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1591_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_1_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5409,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5135_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1492,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_434_I,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5014,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_2_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1472,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1588,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1481,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_CM8I(17),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1588,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_2_36x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4349,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_CM8I(36),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5414,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_2_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1502_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_2_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4977_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_3_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4375_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1429,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_589);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_4_36x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1084,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1044,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_590);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_cm8i_3x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5067,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5411,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1438,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_5303,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_411_I,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_n_23x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1527,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_691_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_o12_n_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1439,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1413,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0(38),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_674_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_x2_0_54x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_440_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_21_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1025,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_4376,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1077,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_21(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(0),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_1x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(1),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_2x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(2),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_3x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(3),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(4),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(5),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(6),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(7),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_8x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(8),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_9x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(9),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(10),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_11x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(11),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_12x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(12),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_13x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(13),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_14x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(14),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_15x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(15),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_16x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(16),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(17),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_18x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(18),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_19x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(19),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_20x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(20),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_21x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(21),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_22x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(22),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_23x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(23),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_24x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(24),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_25x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(25),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_26x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(26),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_27x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(27),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_28x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(28),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_29x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(29),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_30x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(30),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_31x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(31),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_32x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(32),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_33x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(33),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_34x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(34),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_35x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(35),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_36x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(36),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_37x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(37),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_38x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(38),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_39x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(39),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_40x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(40),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_41x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(41),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_42x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(42),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_43x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(43),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_44x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(44),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(45),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_46x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(46),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_47x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(47),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_48x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(48),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_49x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(49),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_50x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(50),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_51x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(51),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_52x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(52),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_53x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(53),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_54x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(54),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_55x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(55),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_56x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(56),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_57x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(57),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_58x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(58),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_59x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(59),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_60x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(60),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_61x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(61),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_62x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(62),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_63x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(63),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_64x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(64),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_65x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(65),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_66x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(66),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_67x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(67),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_68x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(68),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_69x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(69),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_70x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(70),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_71x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(71),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_72x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(72),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_73x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(73),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_74x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(74),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_75x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(75),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_76x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(76),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_77x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(77),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_78x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(78),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_79x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(79),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(80),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(81),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_82x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(82),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_83x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(83),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_84x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(84),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_85x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(85),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_86x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(86),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_87x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(87),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_88x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(88),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_89x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(89),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_90x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(90),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_91x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(91),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_92x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(92),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_93x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(93),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_94x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(94),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_95x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(95),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_96x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(96),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_97x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(97),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_98x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(98),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_99x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(99),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_100x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(100),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_101x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(101),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_102x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(102),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_103x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(103),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_104x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(104),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_105x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(105),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_106x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(106),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_107x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(107),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_108x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(108),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_109x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(109),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_110x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(110),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_111x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(111),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_112x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(112),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_113x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(113),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_114x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(114),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_115x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(115),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_116x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(116),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(116));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_117x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(117),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_118x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(118),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_119x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(119),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_120x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(120),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_121x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(121),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_122x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(122),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_123x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(123),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_124x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(124),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_125x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(125),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_126x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(126),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_127x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(127),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_128x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(128),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_129x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(129),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_130x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(130),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_131x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(131),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_132x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(132),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_133x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(133),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_134x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(134),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_135x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(135),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_136x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(136),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_137x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(137),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_138x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(138),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_139x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(139),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_140x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(140),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_141x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(141),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_142x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(142),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_143x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(143),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_144x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(144),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_145x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(145),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_146x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(146),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_147x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(147),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_148x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(148),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_149x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(149),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_150x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(150),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_151x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(151),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_152x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(152),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_153x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(153),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_154x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(154),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_155x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(155),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_156x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(156),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_157x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(157),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_158x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(158),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_159x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(159),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_160x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(160),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_161x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(161),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_162x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(162),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_163x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(163),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_164x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(164),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_165x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(165),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_166x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(166),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_167x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(167),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_168x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(168),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_169x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(169),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_170x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(170),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_171x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(171),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_172x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(172),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_173x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(173),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(173));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_174x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(174));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_175x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(175));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_176x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(176));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_177x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC_0(54),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(177));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_178x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(53),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(178));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_179x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(52),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(179));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_180x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(51),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(180));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_181x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(50),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(181));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_182x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(49),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(182));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_183x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(48),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(183));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_184x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(47),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(184));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_185x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(46),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(185));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_186x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(45),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(186));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_187x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(44),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(187));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_188x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(43),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(188));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_189x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(42),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(189));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_190x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(41),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(190));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_191x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(40),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_1,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(191));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_192x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(39),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(192));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_193x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(38),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(193));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_194x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(37),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(194));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_195x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(36),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(195));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_196x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(35),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(196));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_197x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(34),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(197));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_198x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(33),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(198));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_199x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(32),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(199));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_200x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(31),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(200));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_201x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(30),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(201));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_202x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(29),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(202));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_203x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(28),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(203));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_204x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(27),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(204));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_205x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(26),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(205));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_206x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(25),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(206));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_207x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(24),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(207));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_208x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(23),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(208));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_209x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(22),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(209));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_210x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(21),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(210));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_211x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(20),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(211));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_212x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(19),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(212));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_213x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(18),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(213));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_214x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(17),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(214));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_215x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(16),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(215));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_216x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(15),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(216));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_217x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(14),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(217));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_218x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(13),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(218));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_219x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(12),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(219));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_220x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(11),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(220));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_221x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(10),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(221));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_222x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(9),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(222));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_223x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(8),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(223));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_224x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(7),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(224));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_225x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(6),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(225));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_226x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(5),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(226));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_227x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(4),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(227));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_228x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(3),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(228));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_229x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(229));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_230x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(230));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_231x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(231));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_232x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(232),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_233x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(233),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_234x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(234),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_235x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(235),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_236x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(236),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_237x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(237),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_238x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(238),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_239x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(239),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_240x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(240),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_241x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(241),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_242x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(242),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_243x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(243),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_244x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(244),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_245x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(245),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_246x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(246),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_247x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(247),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_248x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(248),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_249x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(249),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_250x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(250),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_251x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(251),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_252x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(252),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_253x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(253),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_254x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(254),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_255x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(255),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_256x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(256),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_257x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(257),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_258x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49(258),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(258));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_259x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(0),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_2,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(259));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_260x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(1),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(260));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_261x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(2),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(261));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_262x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(3),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(262));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_263x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(4),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(263));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_264x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(5),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(264));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_265x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(6),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(265));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_266x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(7),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(266));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_267x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(8),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(267));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_268x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(9),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_3,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(268));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_269x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(10),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(269));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_270x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(11),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(270));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_271x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(12),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(271));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_272x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(13),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(272));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_273x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(14),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(273));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_274x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(15),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(274));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_275x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(16),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(275));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_276x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(17),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(276));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_277x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(18),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_4,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(277));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_278x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(19),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(278));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_279x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(20),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(279));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_280x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(21),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(280));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_281x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(22),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(281));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_282x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(23),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(282));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_283x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(24),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(283));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_284x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(25),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(284));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_285x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(26),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(285));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_286x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(27),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_5,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(286));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_287x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(28),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(287));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_288x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(29),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(288));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_289x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(30),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(289));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_290x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(31),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(290));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_291x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(32),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(291));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_292x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(33),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(292));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_293x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(34),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(293));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_294x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(35),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(294));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_295x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(36),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_6,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(295));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_296x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(37),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(296));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_297x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(38),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(297));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_298x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(39),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(298));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_299x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(40),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(299));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_300x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(41),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(300));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_301x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(42),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(301));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_302x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(43),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(302));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_303x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(44),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(303));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_304x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(45),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_7,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(304));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_305x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(46),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(305));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_306x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(47),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(306));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_307x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(48),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(307));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_308x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(49),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(308));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_309x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(50),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(309));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_310x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(51),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(310));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_311x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(52),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(311));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_312x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(53),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(312));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_313x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(54),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_8,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(313));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_314x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(55),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(314));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_315x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(57),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(315));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_316x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_50(316),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_317x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(58),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(317));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_318x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(59),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(318));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_319x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(60),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(319));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_320x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(61),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(320));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_321x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(62),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(321));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_322x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(63),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_9,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(322));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_323x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(64),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(323));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_324x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(65),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(324));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_325x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(66),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(325));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_326x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(67),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(326));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_327x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(68),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(327));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_328x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(69),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(328));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_329x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(70),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(329));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_330x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(71),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(330));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_331x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(72),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_10,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(331));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_332x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(73),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(332));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_333x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(74),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(333));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_334x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(75),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(334));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_335x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(76),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(335));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_336x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(77),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(336));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_337x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(78),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(337));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_338x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(79),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(338));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_339x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(80),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(339));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_340x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(81),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_11,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(340));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_341x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(82),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(341));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_342x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(83),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(342));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_343x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(84),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(343));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_344x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(85),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(344));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_345x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(86),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(345));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_346x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(87),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(346));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_347x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(88),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(347));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_348x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(89),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(348));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_349x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(90),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_12,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(349));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_350x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(91),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(350));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_351x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(92),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(351));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_352x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(93),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(352));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_353x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(94),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(353));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_354x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(95),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(354));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_355x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(96),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(355));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_356x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(97),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(356));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_357x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(98),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(357));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_358x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(99),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_13,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(358));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_359x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(100),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(359));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_360x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(101),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(360));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_361x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(102),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(361));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_362x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(103),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(362));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_363x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(104),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(363));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_364x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(105),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(364));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_365x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(106),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(365));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_366x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(107),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(366));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_367x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(108),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_14,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(367));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_368x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(109),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(368));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_369x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(110),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(369));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_370x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(111),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_371x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(112),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(371));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_372x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(113),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(372));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_373x: DFE1B port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0),
      E => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(373));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_374x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(374),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_375x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(375),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_376x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_DIVMULTV(0),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_377x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_0x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(0),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_1x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(1),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_2x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(2),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_3x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(3),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(4),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(5),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(6),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(7),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_8x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(8),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_9x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(9),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(10),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_11x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(11),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_12x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(12),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_13x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(13),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_14x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(14),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_15x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(15),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_16x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(16),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(17),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_18x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(18),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_19x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(19),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_20x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(20),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_21x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(21),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_22x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(22),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_23x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(23),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_24x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(24),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_25x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(25),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_26x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(26),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_27x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(27),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_28x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(28),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_29x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(29),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_30x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(30),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_31x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(31),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_32x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(32),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_33x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(33),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_34x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(34),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_35x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(35),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_36x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(36),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_37x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(37),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_38x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(38),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_39x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(39),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_40x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(40),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_41x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(41),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_42x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(42),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_43x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(43),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_44x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(44),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(45),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_46x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(46),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_47x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(47),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_48x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(48),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_49x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(49),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_50x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(50),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_51x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(51),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_52x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(52),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_53x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(53),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_54x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(54),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_55x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(55),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_56x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(56),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_57x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(57),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_58x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(58),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_59x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(59),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_61x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(61),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(81),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_90x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(90),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(90));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_103x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(103),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(103));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_105x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(105),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(105));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_107x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(107),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(107));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_111x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(111),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(111));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_0_25x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(25),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0_0_52x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(52),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_1_54x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(54),
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_232x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(232));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_233x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(233));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_234x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(234));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_235x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(235));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_236x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(236));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_237x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(237));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_238x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(238));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_239x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(239));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_240x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(240));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_241x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(241));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_242x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(242));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_243x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(243));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_i_244x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_I(244));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_74,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_73,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_72,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_68,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_66,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_65,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_64,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_63,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_12x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_62,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_13x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_61,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_14x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_60,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_15x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_59,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_16x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_58,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_18x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_56,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_19x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_55,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_20x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_54,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_21x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_22x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_52,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_23x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_51,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_24x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_50,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_25x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_49,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_26x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_48,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_27x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_47,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_28x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_46,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_29x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_45,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_30x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_44,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_31x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_43,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_32x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_42,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_33x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_41,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_34x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_40,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_35x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_39,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_36x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_38,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_38x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_123,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_39x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_122,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_40x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_121,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_41x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_120,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_42x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_43x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_118,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_44x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_46x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_115,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_47x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_114,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_48x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_49x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_112,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_50x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_111,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_51x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_110,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_52x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_53x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_108,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_54x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_107,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_55x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_106,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_56x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_105,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_57x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_104,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_58x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_103,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_59x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_102,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_60x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_101,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_61x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_100,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_62x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_99,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_63x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_98,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_64x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_97,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(64));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_65x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_96,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_66x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_95,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(66));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_67x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_94,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(67));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_68x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_93,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_70x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_91,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(70));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_71x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_90,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_73x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_88,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(73));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_74x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_87,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_75x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_89,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(72));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_76x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_85,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(76));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_77x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_84,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_78x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_83,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_79x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_82,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_82x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_79,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_83x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_78,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_84x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_77,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_85x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_76,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_73,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_68,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_16x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_58,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_11(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_9(18),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_10(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(24),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_646,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(24),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_26x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_48,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_28x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_46,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_29x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_45,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_30x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_44,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_31x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_43,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_32x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_42,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_33x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_41,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_34x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_40,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_36x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_38,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(38),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(37),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_123);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(39),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_674_N,
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_122);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_559,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(40),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(39),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_121);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(40),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_120);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(42),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(41),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(43),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(42),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_118);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(44),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(43),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_4_N(44),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(46),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(46),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1500,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(46),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0(45),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_115);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_21(47),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_114);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(48),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N(47),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(48),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_112);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(50),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_14_N(49),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_111);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(51),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_9_N(50),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_110);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(51),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(53),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19_N(52),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_108);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_107);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_106);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_105);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(57),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(57),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_24_N(56),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_23_N(56),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_104);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(58),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_103);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(59),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(58),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_102);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(60),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(60),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(60),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21(59),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(60),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N(59),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_101);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(61),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(61),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_20_N(60),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(61),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_19_N(60),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_100);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(62),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(61),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_99);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_63x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(63),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(63),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(63),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_6(62),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(63),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5_N(62),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_98);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_64x: OR2A port map (
      A => rst,
      B => GRLFPC2_0_COMB_UN10_IUEXEC,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_97);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_65x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_2_0(65),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(65),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_96);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_66x: AND4B port map (
      A => GRLFPC2_0_COMB_UN10_IUEXEC,
      B => GRLFPC2_0_COMB_UN4_LOCK,
      C => HOLDN_1,
      D => GRLFPC2_0_RS2_0_SQMUXA,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_95);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_67x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(67),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(67),
      D3 => NN_4,
      S00 => NN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      S11 => GRLFPC2_0_FPI_START,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_94);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_68x: OR2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_93);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_70x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_91);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_71x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_FPI_START,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(71),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_90);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_72x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_89);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_73x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN4_NOTRESETORUNIMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_88);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_74x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(62),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_87);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_76x: OR3C port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_TEMP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(61),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_85);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_77x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14_2(77),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_84);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_78x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2051,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_83);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_79x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2040,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_SN_N_19,
      S01 => NN_4,
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_82);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_80x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2049,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_81x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2048,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_82x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2047,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_79);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_83x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2046,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_78);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_84x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2025,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2035,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(84),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(84),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_SN_N_19,
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_77);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_85x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(85),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2034,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_SN_N_19,
      S01 => NN_4,
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_76);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_42x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_44x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_48x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_52x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_65x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_96,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_0_65x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_96,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_0_80x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2049,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_0_0_81x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2048,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2052_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_1_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_38x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_39x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_40x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_42x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_43x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_44x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_45x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_46x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_48x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_50x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_51x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_53x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_57x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_60x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_61x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_63x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_65x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_67x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(67));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_71x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_84x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_0_cm8i_85x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2024_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_CM8I(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N(0),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_74);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_678,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(1),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(1),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_73);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(2),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_72);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(3),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N(3),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_19(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_18_N(6),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_68);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_678,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(8),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_66);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_65);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_464,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(10),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(10),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_64);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_22_N(11),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(11),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_21_N(11),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_63);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(12),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_5_N(12),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_62);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_18(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_17_N(13),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_61);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_1(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(14),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_N(14),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_60);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(15),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_3(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(15),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(15),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_59);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_464,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(16),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2_N(10),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_58);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(17),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_10_N(17),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_19,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_21(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(19),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_20_N(19),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_55);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(20),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_54);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(22),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_646,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(22),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_691_N,
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_52);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_2(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(23),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_691_N,
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_13,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_50);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(25),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_11_N(25),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_49);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_7(26),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(26),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_N(26),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_48);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_47);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_5(28),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(28),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_4_N(28),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1194,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(29),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_3_N(29),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_44);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_42);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_17(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(33),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_16_N(33),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_13(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(34),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_12_N(34),
      S10 => NN_2,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_40);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(35),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(35),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(36),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_38);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_42x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_68,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_31x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_43,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_36x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_38,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_0_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_0_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_0_1_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1_3_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_1_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_0x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_1x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_2x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_3x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_6x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_8x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_10x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_11x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_12x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_13x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_14x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_15x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_16x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_17x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_19x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_22x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_23x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_25x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_26x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_28x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_29x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_33x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_1_cm8i_34x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_68,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_31x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_43,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_42x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_2_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_3_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_4_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_70,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_17x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_57,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_45x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_5_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_6_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_67_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_7_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_8_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_9_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_69_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_80x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_81_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_81x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_80_0,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_10_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_79x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(79),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_83x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(83),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_11_85x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(85),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_12_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_12_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_12_82x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(82),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_12_84x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(84),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_13_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_13_78x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(78),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_14_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_141,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_1x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_140,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_2x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_139,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_3x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_138,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_4x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_5x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_136,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_6x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_135,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_7x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_134,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_8x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_9x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_132,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_11x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_130,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_12x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_129,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_13x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_128,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_14x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_127,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_15x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_126,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_16x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_125,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN58_SCTRL_NEW,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_2,
      S00 => cpi_d_inst(11),
      S01 => cpi_d_inst(9),
      S10 => cpi_d_inst(12),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_141);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_1x: AND4A port map (
      A => cpi_d_inst(12),
      B => cpi_d_inst(11),
      C => cpi_d_inst(7),
      D => cpi_d_inst(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_140);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_2x: AND4B port map (
      A => cpi_d_inst(12),
      B => cpi_d_inst(7),
      C => cpi_d_inst(11),
      D => cpi_d_inst(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_139);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_138);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_4x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(4),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_5x: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_136);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_6x: AND3B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_10(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_135);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_10(10),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_134);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_132);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_10(10),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(11),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_130);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3(0),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_129);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_13x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_AREGSIGN_SEL_INV_1,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(13),
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(13),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPRF_DOUT1_M(63),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_M(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_128);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(14),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_127);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_15x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(15),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_126);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(16),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_125);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_0_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_0_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_0_0_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_1_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_cm8i_11x: CM8INV port map (
      A => cpi_d_inst(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_cm8i_13x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_cm8i_14x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_cm8i_15x: CM8INV port map (
      A => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_1_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_1_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_1_0_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_2_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_2_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_3_10x: DF1 port map (
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
      CLK => clk,
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_3_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_4_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_5_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_6_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_7_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_8_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_9_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_10_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_11_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_12_11x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_0(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_m_12x: AND3A port map (
      A => GRLFPC2_0_FPI_LDOP_2,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_M_0_0(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_M(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_m_0_0_12x: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN2_SIGTAF38_37,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_M_0_0(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2416,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2535,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2476,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2476,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2414,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2533,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2413,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2532,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2473,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2473,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2531,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2412,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2412,
      S00 => N_7988,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2411,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2530,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2410,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2529,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2409,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2528,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(7),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2408,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2527,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(8),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2407,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2526,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2467,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2467,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2406,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2525,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(10),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2405,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2524,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(11),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2404,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2523,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2403,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2522,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2402,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2521,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2401,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2520,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2400,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2519,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(16),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2399,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2518,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2398,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2517,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(18),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2397,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2516,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2396,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2515,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(20),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2395,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2514,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(21),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2394,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2513,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(22),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2393,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2512,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2392,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2511,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(24),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2391,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2510,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2390,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2509,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(26),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2389,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2508,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(27),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2388,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2507,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(28),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2387,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2506,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2386,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2505,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(30),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2385,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2504,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2503,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2384,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2384,
      S00 => N_7988,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2502,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2383,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2383,
      S00 => N_7988,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2382,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2501,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2381,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2500,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2380,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2499,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2379,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2498,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2378,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2497,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2377,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2496,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2376,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2495,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2375,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2494,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2374,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2493,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2373,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2492,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2372,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2491,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2490,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2370,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2489,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2369,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2488,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2368,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2487,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2367,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2486,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2366,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2485,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2365,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2484,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2364,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2483,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2363,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2482,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(53),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2362,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2481,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(54),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2361,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2480,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(55),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2925,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2925,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(58),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2924,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2924,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(59),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2923,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(60),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2922,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(61),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2921,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(62),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_63x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2920,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(63),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_64x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2919,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(64),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(64));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_65x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2918,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(65),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_66x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2917,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(66),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(66));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_67x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2916,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(67),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(67));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_68x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2915,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(68),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_69x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2914,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(69),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(69));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_70x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2913,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(70),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(70));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_71x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2912,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(71),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_72x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2911,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(72),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(72));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_73x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2910,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(73),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(73));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_74x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2909,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(74),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_75x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2908,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(75),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(75));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_76x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2907,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(76),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(76));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_77x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2906,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(77),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_78x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2905,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(78),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_79x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2904,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(79),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_80x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2903,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(80),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_81x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2902,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(81),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_82x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2901,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(82),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_83x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2900,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_0(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(83),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_84x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2899,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(84),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_85x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2898,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(85),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_86x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2897,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(86),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(86));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_87x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2896,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(87),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(87));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_88x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2895,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(88),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(88));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_89x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2894,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(89),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(89));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_90x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2893,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(90),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(90));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_91x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2892,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(91),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(91));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_92x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2891,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(92),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(92));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_93x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2890,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(93),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(93));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_94x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2889,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(94),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(94));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_95x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2888,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2888,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(95),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(95));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_96x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2887,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2887,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(96),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(96));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_97x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2886,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2886,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(97),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(97));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_98x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2885,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(98),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(98));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_99x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2884,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2884,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(99),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(99));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_100x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2883,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2883,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(100),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(100));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_101x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2882,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2882,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(101),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_0(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(101));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_102x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2881,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2881,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(102),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(102));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_103x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2880,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2880,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(103),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(103));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_104x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2879,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2879,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(104),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(104));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_105x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2878,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2878,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(105),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(105));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_106x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2877,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2877,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(106),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(106));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_107x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2876,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2876,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(107),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(107));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_108x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2875,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2875,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(108),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(108));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_109x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2874,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2874,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(109),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(109));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_110x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2873,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2873,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(110),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(110));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_111x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2872,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2872,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(111),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(111));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_112x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2871,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2871,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(112),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(112));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_113x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2870,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2870,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(113),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(113));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_114x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2869,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(114));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_115x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2868,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2868,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(115));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_116x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(116),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(116));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_117x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(117));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_118x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(118));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_119x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
      D1 => GRLFPC2_0_FPO_FRAC(54),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(119));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_120x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
      D1 => GRLFPC2_0_FPO_FRAC(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(120));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_121x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
      D1 => GRLFPC2_0_FPO_FRAC(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(121));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_122x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
      D1 => GRLFPC2_0_FPO_FRAC(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(122));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_123x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
      D1 => GRLFPC2_0_FPO_FRAC(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(123));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_124x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
      D1 => GRLFPC2_0_FPO_FRAC(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(124));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_125x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
      D1 => GRLFPC2_0_FPO_FRAC(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(125));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_126x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
      D1 => GRLFPC2_0_FPO_FRAC(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(126));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_127x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
      D1 => GRLFPC2_0_FPO_FRAC(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(127));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_128x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
      D1 => GRLFPC2_0_FPO_FRAC(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(128));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_129x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
      D1 => GRLFPC2_0_FPO_FRAC(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(129));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_130x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
      D1 => GRLFPC2_0_FPO_FRAC(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(130));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_131x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
      D1 => GRLFPC2_0_FPO_FRAC(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(131));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_132x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
      D1 => GRLFPC2_0_FPO_FRAC(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(132));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_133x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
      D1 => GRLFPC2_0_FPO_FRAC(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(133));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_134x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
      D1 => GRLFPC2_0_FPO_FRAC(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(134));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_135x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
      D1 => GRLFPC2_0_FPO_FRAC(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(135));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_136x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
      D1 => GRLFPC2_0_FPO_FRAC(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(136));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_137x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
      D1 => GRLFPC2_0_FPO_FRAC(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(137));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_138x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
      D1 => GRLFPC2_0_FPO_FRAC(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(138));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_139x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
      D1 => GRLFPC2_0_FPO_FRAC(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(139));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_140x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
      D1 => GRLFPC2_0_FPO_FRAC(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(140));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_141x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3110,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3110,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN8_INFORCREGSN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(141),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(141));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_142x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3109,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14(142),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(142));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_143x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
      D1 => GRLFPC2_0_FPO_FRAC(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(143));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_144x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
      D1 => GRLFPC2_0_FPO_FRAC(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(144));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_145x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
      D1 => GRLFPC2_0_FPO_FRAC(28),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(145));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_146x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
      D1 => GRLFPC2_0_FPO_FRAC(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(146));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_147x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
      D1 => GRLFPC2_0_FPO_FRAC(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(147));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_148x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
      D1 => GRLFPC2_0_FPO_FRAC(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(148));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_149x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
      D1 => GRLFPC2_0_FPO_FRAC(24),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(149));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_150x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
      D1 => GRLFPC2_0_FPO_FRAC(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(150));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_151x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
      D1 => GRLFPC2_0_FPO_FRAC(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(151));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_152x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
      D1 => GRLFPC2_0_FPO_FRAC(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(152));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_153x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
      D1 => GRLFPC2_0_FPO_FRAC(20),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(153));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_154x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
      D1 => GRLFPC2_0_FPO_FRAC(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(154));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_155x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
      D1 => GRLFPC2_0_FPO_FRAC(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(155));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_156x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
      D1 => GRLFPC2_0_FPO_FRAC(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(156));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_157x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
      D1 => GRLFPC2_0_FPO_FRAC(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(157));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_158x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
      D1 => GRLFPC2_0_FPO_FRAC(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(158));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_159x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
      D1 => GRLFPC2_0_FPO_FRAC(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(159));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_160x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
      D1 => GRLFPC2_0_FPO_FRAC(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(160));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_161x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
      D1 => GRLFPC2_0_FPO_FRAC(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(161));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_162x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
      D1 => GRLFPC2_0_FPO_FRAC(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(162));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_163x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
      D1 => GRLFPC2_0_FPO_FRAC(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(163));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_164x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
      D1 => GRLFPC2_0_FPO_FRAC(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(164));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_165x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
      D1 => GRLFPC2_0_FPO_FRAC(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(165));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_166x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
      D1 => GRLFPC2_0_FPO_FRAC(7),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(166));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_167x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
      D1 => GRLFPC2_0_FPO_FRAC(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(167));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_168x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
      D1 => GRLFPC2_0_FPO_FRAC(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(168));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_169x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
      D1 => GRLFPC2_0_FPO_FRAC(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(169));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_170x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
      D1 => GRLFPC2_0_FPO_FRAC(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(170));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_171x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3080,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3080,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_172x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3079,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_QUOBITS(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3079,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(172),
      S11 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(172));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_173x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(173),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(173));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_234x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      D1 => GRLFPC2_0_OP2(62),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3219,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(234),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(234));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_235x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      D1 => GRLFPC2_0_OP2(61),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3218,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(235),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(235));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_236x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      D1 => GRLFPC2_0_OP2(60),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3217,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(236),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(236));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_237x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D1 => GRLFPC2_0_OP2(59),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3206,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3216,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(237),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(237));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_238x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      D1 => GRLFPC2_0_OP2(58),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3205,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3215,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(238),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(238));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_239x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D1 => GRLFPC2_0_OP2(57),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3204,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3214,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(239),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(239));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_240x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D1 => GRLFPC2_0_OP2(56),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3203,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3213,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(240),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(240));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_241x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D1 => GRLFPC2_0_OP2(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3202,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3212,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(241),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(241));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_242x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      D1 => GRLFPC2_0_OP2(54),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3201,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3211,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(242),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(242));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_243x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      D1 => GRLFPC2_0_OP2(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3200,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3210,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(243),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(243));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_244x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      D1 => GRLFPC2_0_OP2(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3199,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3209,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(244),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(244));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_245x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3020,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3006,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(245));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_246x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3019,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3005,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(246));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_247x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3046,
      D1 => NN_2,
      D2 => GRLFPC2_0_OP1(62),
      D3 => NN_2,
      S00 => GRLFPC2_0_FPI_LDOP_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4(11),
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(247));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_248x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3045,
      D1 => NN_2,
      D2 => GRLFPC2_0_OP1(61),
      D3 => NN_2,
      S00 => GRLFPC2_0_FPI_LDOP_2,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(248));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_249x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3016,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3002,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3031,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3031,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(249));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_250x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3015,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3001,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3030,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3030,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(250));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_251x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3014,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3000,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3029,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3029,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(251));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_252x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3013,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2999,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3028,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3028,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(252));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_253x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3012,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2998,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3027,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3027,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(253));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_254x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3011,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2997,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3026,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3026,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(254));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_255x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3010,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2996,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3025,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3025,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(255));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_256x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3009,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2995,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3024,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3024,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(256));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_257x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3008,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2994,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3023,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3023,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_FPI_LDOP_3,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(257));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_374x: OR3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN86_DIVMULTV_N,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN111_DIVMULTV,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0(374),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(374));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_375x: OR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1(375),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0(375),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2120);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      D1 => GRLFPC2_0_FPO_FRAC(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2118);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_3x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(54),
      D1 => GRLFPC2_0_FPO_FRAC(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2117);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_26x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(31),
      D1 => GRLFPC2_0_FPO_FRAC(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2094);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_27x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(30),
      D1 => GRLFPC2_0_FPO_FRAC(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2093);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_28x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(29),
      D1 => GRLFPC2_0_FPO_FRAC(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2092);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_29x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(28),
      D1 => GRLFPC2_0_FPO_FRAC(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2091);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_30x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(27),
      D1 => GRLFPC2_0_FPO_FRAC(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2090);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_31x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(26),
      D1 => GRLFPC2_0_FPO_FRAC(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2089);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_32x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(25),
      D1 => GRLFPC2_0_FPO_FRAC(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2088);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_33x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(24),
      D1 => GRLFPC2_0_FPO_FRAC(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2087);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_34x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(23),
      D1 => GRLFPC2_0_FPO_FRAC(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2086);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_35x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(22),
      D1 => GRLFPC2_0_FPO_FRAC(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2085);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_36x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(21),
      D1 => GRLFPC2_0_FPO_FRAC(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2084);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_37x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(20),
      D1 => GRLFPC2_0_FPO_FRAC(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2083);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_38x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(19),
      D1 => GRLFPC2_0_FPO_FRAC(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2082);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_39x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(18),
      D1 => GRLFPC2_0_FPO_FRAC(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2081);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_40x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(17),
      D1 => GRLFPC2_0_FPO_FRAC(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2080);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_41x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(16),
      D1 => GRLFPC2_0_FPO_FRAC(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2079);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_42x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(15),
      D1 => GRLFPC2_0_FPO_FRAC(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2078);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_43x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(14),
      D1 => GRLFPC2_0_FPO_FRAC(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2077);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_44x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(13),
      D1 => GRLFPC2_0_FPO_FRAC(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2076);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_45x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(12),
      D1 => GRLFPC2_0_FPO_FRAC(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2075);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_46x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(11),
      D1 => GRLFPC2_0_FPO_FRAC(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2074);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_47x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(10),
      D1 => GRLFPC2_0_FPO_FRAC(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2073);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_48x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(9),
      D1 => GRLFPC2_0_FPO_FRAC(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2072);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_49x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(8),
      D1 => GRLFPC2_0_FPO_FRAC(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2071);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_50x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(7),
      D1 => GRLFPC2_0_FPO_FRAC(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2070);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_51x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(6),
      D1 => GRLFPC2_0_FPO_FRAC(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2069);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_52x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(5),
      D1 => GRLFPC2_0_FPO_FRAC(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2068);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_53x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(4),
      D1 => GRLFPC2_0_FPO_FRAC(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2067);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_54x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2066);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2065);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2064);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_57x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2063);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_58x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2746);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_59x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      D1 => GRLFPC2_0_FPO_FRAC(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2745);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      D1 => GRLFPC2_0_FPO_FRAC(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2744);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_84x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(31),
      D1 => GRLFPC2_0_FPO_FRAC(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2720);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_85x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(30),
      D1 => GRLFPC2_0_FPO_FRAC(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2719);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_86x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(29),
      D1 => GRLFPC2_0_FPO_FRAC(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2718);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_87x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(28),
      D1 => GRLFPC2_0_FPO_FRAC(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2717);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_88x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(27),
      D1 => GRLFPC2_0_FPO_FRAC(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2716);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_89x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(26),
      D1 => GRLFPC2_0_FPO_FRAC(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2715);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_90x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(25),
      D1 => GRLFPC2_0_FPO_FRAC(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2714);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_91x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(24),
      D1 => GRLFPC2_0_FPO_FRAC(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2713);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_92x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(23),
      D1 => GRLFPC2_0_FPO_FRAC(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2712);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_93x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(22),
      D1 => GRLFPC2_0_FPO_FRAC(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2711);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_94x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(21),
      D1 => GRLFPC2_0_FPO_FRAC(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2710);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_95x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(20),
      D1 => GRLFPC2_0_FPO_FRAC(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2709);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_96x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(19),
      D1 => GRLFPC2_0_FPO_FRAC(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2708);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_97x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(18),
      D1 => GRLFPC2_0_FPO_FRAC(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2707);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_98x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(17),
      D1 => GRLFPC2_0_FPO_FRAC(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2706);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_99x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(16),
      D1 => GRLFPC2_0_FPO_FRAC(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2705);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_100x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(15),
      D1 => GRLFPC2_0_FPO_FRAC(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2704);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_101x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(14),
      D1 => GRLFPC2_0_FPO_FRAC(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2703);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_102x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(13),
      D1 => GRLFPC2_0_FPO_FRAC(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2702);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_103x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(12),
      D1 => GRLFPC2_0_FPO_FRAC(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2701);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_104x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(11),
      D1 => GRLFPC2_0_FPO_FRAC(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2700);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_105x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(10),
      D1 => GRLFPC2_0_FPO_FRAC(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2699);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_106x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(9),
      D1 => GRLFPC2_0_FPO_FRAC(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2698);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_107x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(8),
      D1 => GRLFPC2_0_FPO_FRAC(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2697);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_108x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(7),
      D1 => GRLFPC2_0_FPO_FRAC(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2696);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_109x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(6),
      D1 => GRLFPC2_0_FPO_FRAC(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2695);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_110x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(5),
      D1 => GRLFPC2_0_FPO_FRAC(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2694);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_111x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2693);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_112x: CM8 port map (
      D0 => GRLFPC2_0_FPO_FRAC(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2692);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_113x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2691);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_114x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2690);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_115x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2689);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_141x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
      D1 => GRLFPC2_0_FPO_FRAC(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3110);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_142x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
      D1 => GRLFPC2_0_FPO_FRAC(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3109);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_171x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I(171),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3080);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_172x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I(172),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3079);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_237x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      D1 => GRLFPC2_0_OP2(62),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3206);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_238x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      D1 => GRLFPC2_0_OP2(61),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3205);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_239x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D1 => GRLFPC2_0_OP2(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3204);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_240x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D1 => GRLFPC2_0_OP2(59),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3203);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_241x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(7),
      D1 => GRLFPC2_0_OP2(58),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3202);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_242x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D1 => GRLFPC2_0_OP2(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3201);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_243x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D1 => GRLFPC2_0_OP2(56),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3200);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_244x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D1 => GRLFPC2_0_OP2(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3199);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_245x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3006);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_246x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3005);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_247x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3004);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_248x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3003);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_249x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3002);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_250x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3001);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_251x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(6),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3000);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_252x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(5),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2999);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_253x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2998);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_254x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2997);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_255x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2996);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_256x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2995);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_257x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2994);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_374x: XOR2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0(374));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_375x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTDIVISORBIT,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I(375),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_cm8i_171x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_cm8i_172x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I(172));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_cm8i_375x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_CM8I(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2178);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2176);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      D1 => GRLFPC2_0_OP2(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      D3 => GRLFPC2_0_OP2(53),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2175);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D1 => GRLFPC2_0_OP2(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D3 => GRLFPC2_0_OP2(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2174);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D1 => GRLFPC2_0_OP2(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D3 => GRLFPC2_0_OP2(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2173);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D1 => GRLFPC2_0_OP2(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D3 => GRLFPC2_0_OP2(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2172);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D1 => GRLFPC2_0_OP2(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D3 => GRLFPC2_0_OP2(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2171);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D1 => GRLFPC2_0_OP2(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D3 => GRLFPC2_0_OP2(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2170);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D1 => GRLFPC2_0_OP2(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D3 => GRLFPC2_0_OP2(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2169);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D1 => GRLFPC2_0_OP2(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D3 => GRLFPC2_0_OP2(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2168);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D1 => GRLFPC2_0_OP2(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D3 => GRLFPC2_0_OP2(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2167);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      D1 => GRLFPC2_0_OP2(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      D3 => GRLFPC2_0_OP2(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2166);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D1 => GRLFPC2_0_OP2(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D3 => GRLFPC2_0_OP2(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2165);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D1 => GRLFPC2_0_OP2(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D3 => GRLFPC2_0_OP2(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2164);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D1 => GRLFPC2_0_OP2(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D3 => GRLFPC2_0_OP2(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2163);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D1 => GRLFPC2_0_OP2(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D3 => GRLFPC2_0_OP2(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2162);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      D1 => GRLFPC2_0_OP2(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(18),
      D3 => GRLFPC2_0_OP2(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2161);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      D1 => GRLFPC2_0_OP2(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(19),
      D3 => GRLFPC2_0_OP2(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2160);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D1 => GRLFPC2_0_OP2(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D3 => GRLFPC2_0_OP2(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2159);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      D1 => GRLFPC2_0_OP2(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(21),
      D3 => GRLFPC2_0_OP2(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2158);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D1 => GRLFPC2_0_OP2(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D3 => GRLFPC2_0_OP2(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2157);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      D1 => rfo2_data2(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(23),
      D3 => GRLFPC2_0_OP2(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2156);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      D1 => rfo2_data2(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      D3 => GRLFPC2_0_OP2(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2155);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D1 => rfo2_data2(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D3 => GRLFPC2_0_OP2(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2154);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2126);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(54),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2125);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_56x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2123);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN7_XZAREGLOADEN,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL_0_0,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      D1 => GRLFPC2_0_OP1(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      D3 => GRLFPC2_0_OP1(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2802);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      D1 => GRLFPC2_0_OP1(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      D3 => GRLFPC2_0_OP1(53),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2801);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_63x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      D1 => GRLFPC2_0_OP1(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      D3 => GRLFPC2_0_OP1(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2800);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_64x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      D1 => GRLFPC2_0_OP1(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      D3 => GRLFPC2_0_OP1(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2799);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_65x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      D1 => GRLFPC2_0_OP1(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      D3 => GRLFPC2_0_OP1(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2798);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_66x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      D1 => GRLFPC2_0_OP1(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      D3 => GRLFPC2_0_OP1(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2797);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_67x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      D1 => GRLFPC2_0_OP1(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      D3 => GRLFPC2_0_OP1(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2796);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_68x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      D1 => GRLFPC2_0_OP1(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      D3 => GRLFPC2_0_OP1(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2795);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_69x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      D1 => GRLFPC2_0_OP1(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      D3 => GRLFPC2_0_OP1(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2794);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_70x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      D1 => GRLFPC2_0_OP1(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      D3 => GRLFPC2_0_OP1(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2793);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_71x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      D1 => GRLFPC2_0_OP1(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      D3 => GRLFPC2_0_OP1(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2792);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_72x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      D1 => GRLFPC2_0_OP1(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      D3 => GRLFPC2_0_OP1(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2791);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_73x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      D1 => GRLFPC2_0_OP1(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      D3 => GRLFPC2_0_OP1(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2790);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_74x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      D1 => GRLFPC2_0_OP1(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      D3 => GRLFPC2_0_OP1(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2789);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_75x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      D1 => GRLFPC2_0_OP1(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      D3 => GRLFPC2_0_OP1(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2788);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_76x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      D1 => GRLFPC2_0_OP1(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      D3 => GRLFPC2_0_OP1(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2787);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_77x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      D1 => GRLFPC2_0_OP1(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      D3 => GRLFPC2_0_OP1(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2786);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_78x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      D1 => GRLFPC2_0_OP1(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      D3 => GRLFPC2_0_OP1(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2785);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_79x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      D1 => GRLFPC2_0_OP1(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      D3 => GRLFPC2_0_OP1(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2784);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_80x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      D1 => GRLFPC2_0_OP1(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      D3 => GRLFPC2_0_OP1(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2783);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_81x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      D1 => rfo2_data1(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      D3 => GRLFPC2_0_OP1(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2782);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_82x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      D1 => rfo2_data1(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      D3 => GRLFPC2_0_OP1(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2781);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_83x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      D1 => rfo2_data1(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      D3 => GRLFPC2_0_OP1(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2780);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_95x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(95),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2768);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_96x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(96),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2767);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_97x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(97),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2766);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_99x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(99),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2764);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_100x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(100),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2763);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_101x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(101),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2762);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_102x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(102),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2761);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_103x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(103),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2760);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_104x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(104),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2759);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_105x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(105),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2758);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_106x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(106),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2757);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_107x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(107),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2756);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_108x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(108),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2755);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_109x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(109),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2754);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_110x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(110),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2753);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_111x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(111),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2752);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_112x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(112),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2751);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_232x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3221);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_233x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3220);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_234x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(10),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3219);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_235x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3218);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_236x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(8),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3217);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_237x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3216);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_238x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(6),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3215);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_239x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(5),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3214);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_240x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3213);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_241x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3212);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_242x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLC(0),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3211);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_243x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3210);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_244x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3209);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_245x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3020);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_246x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3019);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_249x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      D1 => GRLFPC2_0_FPO_EXP(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3016);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_250x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      D1 => GRLFPC2_0_FPO_EXP(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3015);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_251x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      D1 => GRLFPC2_0_FPO_EXP(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3014);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_252x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      D1 => GRLFPC2_0_FPO_EXP(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3013);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_253x: CM8 port map (
      D0 => GRLFPC2_0_FPO_EXP(5),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_15,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3067,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3012);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_254x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      D1 => GRLFPC2_0_FPO_EXP(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3011);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_255x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      D1 => GRLFPC2_0_FPO_EXP(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3010);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_256x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      D1 => GRLFPC2_0_FPO_EXP(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3009);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_257x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      D1 => GRLFPC2_0_FPO_EXP(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3008);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_375x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTDIVISORBIT,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_95x: CM8INV port map (
      A => rfo2_data1(17),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(95));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_96x: CM8INV port map (
      A => rfo2_data1(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(96));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_97x: CM8INV port map (
      A => rfo2_data1(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(97));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_99x: CM8INV port map (
      A => rfo2_data1(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(99));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_100x: CM8INV port map (
      A => rfo2_data1(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(100));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_101x: CM8INV port map (
      A => rfo2_data1(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(101));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_102x: CM8INV port map (
      A => rfo2_data1(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(102));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_103x: CM8INV port map (
      A => rfo2_data1(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(103));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_104x: CM8INV port map (
      A => rfo2_data1(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(104));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_105x: CM8INV port map (
      A => rfo2_data1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(105));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_106x: CM8INV port map (
      A => rfo2_data1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(106));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_107x: CM8INV port map (
      A => rfo2_data1(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(107));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_108x: CM8INV port map (
      A => rfo2_data1(4),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(108));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_109x: CM8INV port map (
      A => rfo2_data1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(109));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_110x: CM8INV port map (
      A => rfo2_data1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(110));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_111x: CM8INV port map (
      A => rfo2_data1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(111));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_cm8i_112x: CM8INV port map (
      A => rfo2_data1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_CM8I(112));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2234);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2233);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2232);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2231);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2230);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2229);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2228);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2226);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2225);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2224);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2223);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2222);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2221);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2220);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2219);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2218);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2217);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2216);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2215);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2214);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2213);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2212);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2211);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2210);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2209);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2208);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(33),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(34),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2206);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(35),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2205);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2204);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(37),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2203);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(38),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2202);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(39),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2201);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(42),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2198);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2194);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2193);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2192);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2191);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2190);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2189);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2188);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2187);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_249x: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      B => GRLFPC2_0_OP1(60),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3031);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_250x: CM8 port map (
      D0 => GRLFPC2_0_OP1(59),
      D1 => GRLFPC2_0_OP1(62),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3030);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_251x: CM8 port map (
      D0 => GRLFPC2_0_OP1(58),
      D1 => GRLFPC2_0_OP1(61),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3029);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_252x: CM8 port map (
      D0 => GRLFPC2_0_OP1(57),
      D1 => GRLFPC2_0_OP1(60),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3028);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_253x: CM8 port map (
      D0 => GRLFPC2_0_OP1(56),
      D1 => GRLFPC2_0_OP1(59),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3027);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_254x: CM8 port map (
      D0 => GRLFPC2_0_OP1(55),
      D1 => GRLFPC2_0_OP1(58),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3026);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_255x: CM8 port map (
      D0 => GRLFPC2_0_OP1(54),
      D1 => GRLFPC2_0_OP1(57),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3025);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_256x: CM8 port map (
      D0 => GRLFPC2_0_OP1(53),
      D1 => GRLFPC2_0_OP1(56),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3024);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_257x: CM8 port map (
      D0 => GRLFPC2_0_OP1(52),
      D1 => GRLFPC2_0_OP1(55),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12(11),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3023);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_58x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2746,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(58),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2925);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_59x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2745,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(59),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2924);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_60x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2744,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2744,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2923);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_61x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2802,
      D1 => GRLFPC2_0_FPO_FRAC(54),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2802,
      D3 => GRLFPC2_0_FPO_FRAC(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2922);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_62x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2801,
      D1 => GRLFPC2_0_FPO_FRAC(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2801,
      D3 => GRLFPC2_0_FPO_FRAC(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2921);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_63x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2800,
      D1 => GRLFPC2_0_FPO_FRAC(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2800,
      D3 => GRLFPC2_0_FPO_FRAC(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2920);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_64x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2799,
      D1 => GRLFPC2_0_FPO_FRAC(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2799,
      D3 => GRLFPC2_0_FPO_FRAC(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2919);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_65x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2798,
      D1 => GRLFPC2_0_FPO_FRAC(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2798,
      D3 => GRLFPC2_0_FPO_FRAC(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2918);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_66x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2797,
      D1 => GRLFPC2_0_FPO_FRAC(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2797,
      D3 => GRLFPC2_0_FPO_FRAC(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2917);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_67x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2796,
      D1 => GRLFPC2_0_FPO_FRAC(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2796,
      D3 => GRLFPC2_0_FPO_FRAC(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2916);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_68x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2795,
      D1 => GRLFPC2_0_FPO_FRAC(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2795,
      D3 => GRLFPC2_0_FPO_FRAC(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2915);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_69x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2794,
      D1 => GRLFPC2_0_FPO_FRAC(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2794,
      D3 => GRLFPC2_0_FPO_FRAC(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2914);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_70x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2793,
      D1 => GRLFPC2_0_FPO_FRAC(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2793,
      D3 => GRLFPC2_0_FPO_FRAC(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2913);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_71x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2792,
      D1 => GRLFPC2_0_FPO_FRAC(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2792,
      D3 => GRLFPC2_0_FPO_FRAC(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2912);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_72x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2791,
      D1 => GRLFPC2_0_FPO_FRAC(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2791,
      D3 => GRLFPC2_0_FPO_FRAC(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2911);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_73x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2790,
      D1 => GRLFPC2_0_FPO_FRAC(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2790,
      D3 => GRLFPC2_0_FPO_FRAC(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2910);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_74x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2789,
      D1 => GRLFPC2_0_FPO_FRAC(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2789,
      D3 => GRLFPC2_0_FPO_FRAC(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2909);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_75x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2788,
      D1 => GRLFPC2_0_FPO_FRAC(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2788,
      D3 => GRLFPC2_0_FPO_FRAC(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2908);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_76x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2787,
      D1 => GRLFPC2_0_FPO_FRAC(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2787,
      D3 => GRLFPC2_0_FPO_FRAC(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2907);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_77x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2786,
      D1 => GRLFPC2_0_FPO_FRAC(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2786,
      D3 => GRLFPC2_0_FPO_FRAC(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2906);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_78x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2785,
      D1 => GRLFPC2_0_FPO_FRAC(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2785,
      D3 => GRLFPC2_0_FPO_FRAC(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2905);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_79x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2784,
      D1 => GRLFPC2_0_FPO_FRAC(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2784,
      D3 => GRLFPC2_0_FPO_FRAC(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2904);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_80x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2783,
      D1 => GRLFPC2_0_FPO_FRAC(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2783,
      D3 => GRLFPC2_0_FPO_FRAC(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2903);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_81x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2782,
      D1 => GRLFPC2_0_FPO_FRAC(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2782,
      D3 => GRLFPC2_0_FPO_FRAC(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2902);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_82x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2781,
      D1 => GRLFPC2_0_FPO_FRAC(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2781,
      D3 => GRLFPC2_0_FPO_FRAC(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2901);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_83x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2780,
      D1 => GRLFPC2_0_FPO_FRAC(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2780,
      D3 => GRLFPC2_0_FPO_FRAC(30),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2900);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_84x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2720,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(84),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2720,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2899);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_85x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2719,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(85),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2719,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_4,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2898);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_86x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2718,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(86),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2718,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2897);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_87x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2717,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(87),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2717,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2896);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_88x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2716,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(88),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2716,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2895);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_89x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2715,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(89),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2715,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2894);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_90x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2714,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(90),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2714,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2893);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_91x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2713,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(91),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2713,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2892);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_92x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2712,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(92),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2712,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2891);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_93x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2711,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(93),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2711,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2890);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_94x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2710,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(94),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2710,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2889);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_95x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2768,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2709,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2888);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_96x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2767,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2708,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2887);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_97x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2766,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2707,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2886);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_98x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2706,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(98),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2706,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2885);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_99x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2764,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2705,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2884);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_100x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2763,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2704,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2883);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_101x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2762,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2703,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2882);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_102x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2761,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2702,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2881);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_103x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2760,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2701,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2880);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_104x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2759,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2700,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2879);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_105x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2758,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2699,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2878);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_106x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2757,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2698,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2877);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_107x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2756,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2697,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2876);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_108x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2755,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2696,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2875);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_109x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2754,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2695,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2874);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_110x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2753,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2694,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2873);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_111x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2752,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2693,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2872);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_112x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2751,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2692,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2871);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_113x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2691,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(113),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2870);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_114x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2690,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2690,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2869);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_115x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2689,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(115),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2868);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_232x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3221,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(232));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_233x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3220,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(233));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_247x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3004,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3004,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3046);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_248x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      D1 => GRLFPC2_0_FPO_EXP(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3003,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3003,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_UN6_EXPBREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3045);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_cm8i_58x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_cm8i_59x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(59));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_cm8i_113x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(113));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_cm8i_115x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_3_CM8I(115));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_3x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2353);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2347);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_0x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2120,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2120,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_5_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2416);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2118,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2118,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2414);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2176,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2117,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2413);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2175,
      D1 => GRLFPC2_0_FPO_FRAC(53),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2175,
      D3 => GRLFPC2_0_FPO_FRAC(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2412);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2174,
      D1 => GRLFPC2_0_FPO_FRAC(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2174,
      D3 => GRLFPC2_0_FPO_FRAC(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2411);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2173,
      D1 => GRLFPC2_0_FPO_FRAC(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2173,
      D3 => GRLFPC2_0_FPO_FRAC(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2410);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2172,
      D1 => GRLFPC2_0_FPO_FRAC(50),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2172,
      D3 => GRLFPC2_0_FPO_FRAC(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2409);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2171,
      D1 => GRLFPC2_0_FPO_FRAC(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2171,
      D3 => GRLFPC2_0_FPO_FRAC(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2408);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2170,
      D1 => GRLFPC2_0_FPO_FRAC(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2170,
      D3 => GRLFPC2_0_FPO_FRAC(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2407);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2169,
      D1 => GRLFPC2_0_FPO_FRAC(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2169,
      D3 => GRLFPC2_0_FPO_FRAC(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2406);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2168,
      D1 => GRLFPC2_0_FPO_FRAC(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2168,
      D3 => GRLFPC2_0_FPO_FRAC(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2405);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2167,
      D1 => GRLFPC2_0_FPO_FRAC(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2167,
      D3 => GRLFPC2_0_FPO_FRAC(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2404);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2166,
      D1 => GRLFPC2_0_FPO_FRAC(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2166,
      D3 => GRLFPC2_0_FPO_FRAC(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2403);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2165,
      D1 => GRLFPC2_0_FPO_FRAC(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2165,
      D3 => GRLFPC2_0_FPO_FRAC(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2402);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2164,
      D1 => GRLFPC2_0_FPO_FRAC(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2164,
      D3 => GRLFPC2_0_FPO_FRAC(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2401);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2163,
      D1 => GRLFPC2_0_FPO_FRAC(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2163,
      D3 => GRLFPC2_0_FPO_FRAC(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2400);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2162,
      D1 => GRLFPC2_0_FPO_FRAC(40),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2162,
      D3 => GRLFPC2_0_FPO_FRAC(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2399);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2161,
      D1 => GRLFPC2_0_FPO_FRAC(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2161,
      D3 => GRLFPC2_0_FPO_FRAC(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2398);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2160,
      D1 => GRLFPC2_0_FPO_FRAC(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2160,
      D3 => GRLFPC2_0_FPO_FRAC(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2397);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2159,
      D1 => GRLFPC2_0_FPO_FRAC(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2159,
      D3 => GRLFPC2_0_FPO_FRAC(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2396);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2158,
      D1 => GRLFPC2_0_FPO_FRAC(36),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2158,
      D3 => GRLFPC2_0_FPO_FRAC(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2395);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2157,
      D1 => GRLFPC2_0_FPO_FRAC(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2157,
      D3 => GRLFPC2_0_FPO_FRAC(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2394);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2156,
      D1 => GRLFPC2_0_FPO_FRAC(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2156,
      D3 => GRLFPC2_0_FPO_FRAC(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2393);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2155,
      D1 => GRLFPC2_0_FPO_FRAC(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2155,
      D3 => GRLFPC2_0_FPO_FRAC(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2392);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2154,
      D1 => GRLFPC2_0_FPO_FRAC(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2154,
      D3 => GRLFPC2_0_FPO_FRAC(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2391);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2094,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2094,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2390);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2093,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2093,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2389);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2092,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2092,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2388);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2091,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2091,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_5,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2387);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2090,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2090,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2386);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2089,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2089,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2385);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2088,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2088,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2384);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2087,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2087,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2383);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2086,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2086,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2382);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2085,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2085,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2381);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2084,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2084,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2380);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2083,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2083,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2379);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2082,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2082,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_6,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2378);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2081,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2081,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2377);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2080,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2080,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2376);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2079,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2079,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2375);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2078,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2078,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2374);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2077,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2077,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2373);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2076,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2076,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2372);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0(45),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2075,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2075,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2074,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2074,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2370);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2073,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2073,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_7,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2369);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2072,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2072,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2368);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2071,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2071,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2367);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2070,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2070,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2366);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2069,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2069,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2365);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2068,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2068,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2364);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2126,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2067,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2363);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2125,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2066,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2362);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_55x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2065,
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2065,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_5_CM8I(55),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2361);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_5_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_5_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_5_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N(57),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_N(56),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2476);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_N(56),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2_N(56),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2475);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(54),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2353,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2353,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2473);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(48),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2347,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2347,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2467);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_57x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(57),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3288,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2419);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(55),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_6_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(55),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2474_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(53),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(52),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2472_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(52),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2471_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(51),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(50),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2470_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(50),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2469_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(49),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(48),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2468_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(47),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(46),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2466_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(46),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2465_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(45),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2464_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(44),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2463_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(43),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2462_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(42),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2461_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(41),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2460_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(40),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2459_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(39),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2458_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(38),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2457_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(37),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(36),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2456_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(36),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2455_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(35),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2454_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(34),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2453_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(33),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2452_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(32),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2451_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(31),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(30),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2450_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(30),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2449_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(29),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(28),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2448_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(28),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(27),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2447_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(27),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(26),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2446_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(26),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2445_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(25),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(24),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2444_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(24),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2443_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(23),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(22),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2442_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(22),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(21),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2441_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(21),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(20),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2440_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(20),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2439_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(19),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(18),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2438_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(18),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2437_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(17),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(16),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2436_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(16),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2435_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(15),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2434_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(14),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2433_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(13),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2432_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(12),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(11),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2431_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(11),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(10),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2430_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(10),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2429_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(9),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(8),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2428_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(8),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(7),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2427_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(7),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2426_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(6),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_5(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2425_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(5),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(4),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2424_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(4),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2423_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(3),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2422_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(2),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2421_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_6_n_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1(1),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2420_N);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(116),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2535);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2534);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2533);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2532);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2531);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2234,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2234,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2530);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2233,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2233,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2529);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2232,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2232,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2528);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2231,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(8),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2231,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2527);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2230,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2230,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2526);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2229,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(10),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2229,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2525);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2228,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2228,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2524);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2523);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2226,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2226,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2522);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2225,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2225,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2521);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2224,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2224,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2520);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2223,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2223,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2519);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2222,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2222,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2518);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2221,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2221,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2517);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2220,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2220,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2516);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2219,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2219,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2515);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2218,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2218,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2514);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2217,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2217,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2513);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2216,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2216,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2512);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2215,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(24),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2215,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2511);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2214,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2214,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2510);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2213,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2213,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2509);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2212,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2212,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2508);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2211,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(28),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2211,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2507);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2210,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2210,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2506);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2209,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2209,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2505);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2208,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2208,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2504);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(32),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2503);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2206,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2206,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2502);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2205,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2205,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2501);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2204,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2204,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2500);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2203,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(36),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2203,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2499);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2202,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2202,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2498);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2201,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2201,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2497);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2496);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2495);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2198,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2198,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2494);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2493);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2492);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(44),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2491);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2194,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2194,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2490);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2193,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2193,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2489);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2192,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2192,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2488);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2191,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(48),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2191,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2487);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2190,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2190,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2486);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2189,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2189,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_10(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2485);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2188,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2188,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2484);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2187,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2187,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2483);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2482);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(54),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2481);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_7_CM8I(55),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2480);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2479);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(173),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(57),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2478);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_7_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_7_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2474_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_4x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2472_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2471_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_6x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2470_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2469_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_8x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2468_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2466_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2465_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2464_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2463_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2462_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2461_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2460_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2459_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_18x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2458_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2457_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_20x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2456_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2455_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_22x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2454_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2453_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_24x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2452_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2451_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_26x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2450_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2449_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_28x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2448_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2447_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_30x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2446_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_31x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2445_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_32x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2444_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_33x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2443_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_34x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2442_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_35x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2441_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_36x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2440_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_37x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2439_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_38x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2438_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_39x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2437_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_40x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2436_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_41x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2435_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_42x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2434_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2433_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_44x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2432_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2431_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_46x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2430_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2429_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_48x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2428_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_49x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2427_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2426_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2425_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2424_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2423_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2422_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_55x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2421_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_141x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(141));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_172x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(172));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_234x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(234));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_235x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(235));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_236x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(236));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_237x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(237));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_238x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(238));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_239x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(239));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_240x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(240));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_241x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(241));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_242x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(242));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_243x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(243));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_cm8i_244x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_CM8I(244));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_d_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2178,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2475,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2475,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S11 => NN_2,
      Y => N_7984);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_d_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2123,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_D_CM8I(56),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2064,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_D_CM8I(56),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S11 => NN_2,
      Y => N_7983);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_d_57x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2419,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2063,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2419,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6,
      S11 => NN_2,
      Y => N_7980);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_d_cm8i_56x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2420_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_D_CM8I(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_s_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      S11 => NN_2,
      Y => N_7988);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_s_57x: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_S_CM8I(57),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      S11 => NN_2,
      Y => N_7979);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_s_cm8i_57x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_S_CM8I(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_1: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_1_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_2: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_3: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_4: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m2_5: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3076_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_1: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_2: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_3: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_4: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_5: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3136_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_1_0: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3268_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_e: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_e_0: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_e_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_e_2: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_e_3: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1_0_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_S,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_CM8I,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN3_PREVENTSWAP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      D3 => NN_2,
      S00 => GRLFPC2_0_FPI_LDOP_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN5_XZBREGLOADEN_1,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_0_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2866_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0_6: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_6: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_cm8i: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_s: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_FPI_LDOP_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_S);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m5: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_0_SQMUXA_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m5_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_0,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_0_SQMUXA_1_0,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLC_1(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3251_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m5_e: AND2B port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3067);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M6_0_CM8I,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_1(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_0: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_0_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_0_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_1: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_2: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_3: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_4: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_5: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_0_0,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2926_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_FPI_LDOP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M6_0_CM8I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_1: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_2: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_3: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_4: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m6_5: AND2A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(7),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2477_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m7: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_S,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m7_0: AND3A port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_1(5),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M4_S,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m8: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m8_0: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m8_1: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m8_2: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m8_3: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m8_4: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2357_0,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2(6),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2536_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10_0: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10_1: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10_2: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10_3: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10_4: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m10_5: AND3 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_8_0,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1(6),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2595_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(2),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(1),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(2),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(4),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(2),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(4),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(3),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(4),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(4),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(6),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(7),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(6),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_6x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_7x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(9),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_9x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(10),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(11),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(12),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(14),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(16),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(19),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_19x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(21),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_21x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_22x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(23),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_23x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_24x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(25),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_25x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(25),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_26x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(27),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_27x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(29),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_29x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(29),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_30x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(31),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_35x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_37x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_39x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(39),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_42x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_43x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_44x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(45),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_45x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(45),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_46x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(47),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_47x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_48x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(49),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_54x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(55),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_10x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_11x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_12x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_14x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_15x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_16x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_5x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(7),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(5),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_6x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(8),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(6),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(7),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(10),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(8),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_9x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_10x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(12),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(10),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_12x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(14),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(12),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_14x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(16),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(14),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_16x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(18),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(16),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_18x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(18),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_20x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(22),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(20),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_21x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(21),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_22x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(24),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(22),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_24x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(26),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(24),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_25x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_26x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(28),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(26),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_28x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(28),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_29x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_30x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(32),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(30),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_31x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(33),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_32x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(34),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(32),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_33x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(35),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(33),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_34x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(36),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(34),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_35x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(37),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(35),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_36x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(38),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(36),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_37x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(37),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_38x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(38),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_39x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_40x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_41x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_42x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(45),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_44x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(45),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_46x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(48),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_47x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(49),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_48x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(50),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(48),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_49x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_51x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(51),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_52x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(52),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_53x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_54x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_55x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_56x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_7x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(7),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_9x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(11),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_19x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_21x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_23x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(23),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_25x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_27x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(27),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_29x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(31),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_43x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_47x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_50x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(50),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_51x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_52x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_53x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(53),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_cm8i_54x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(54),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2_CM8I(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_2x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_6x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_7x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_8x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_10x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_11x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_12x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_13x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(13),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_14x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_15x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_16x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_17x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_18x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_19x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_20x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_22x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_23x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_24x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_26x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_27x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_28x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_4(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_30x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_31x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_32x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_33x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_34x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_35x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_36x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_37x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_38x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_5(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_39x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_40x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_0(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_41x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_42x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_43x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(47),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_44x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(1),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_46x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(3),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_48x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(1),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(5),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_50x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(3),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(54),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_6(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_cm8i_5x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_cm8i_13x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_cm8i_17x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_CM8I(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_n_45x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(45),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N_CM8I(45),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_n_49x: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(53),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_n_cm8i_45x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_N(49),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2_N_CM8I(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_temp: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_temp_0: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_temp_1: AND2 port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0(42),
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_1x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_3x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_4x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_5x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_n_8x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_N(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_aregsign_sel_inv_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_4,
      D2 => NN_4,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN2_SIGTAF38_37,
      S11 => GRLFPC2_0_FPI_LDOP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_AREGSIGN_SEL_INV_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_divmultv_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_DIVMULTV_CM8I(0),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN5_DIVMULTV,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_DIVMULTV(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_divmultv_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_DIVMULTV_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_0x: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_N,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_CM8I(0),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP_N,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_1_0x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN16_NOTPROP,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1_N(1),
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_GEN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_2_0x: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
      D2 => NN_2,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_NOTPROP,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN47_GEN,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_3_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3_CM8I(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_3,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_3_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN2_NOTPROP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_4: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      fci => NN_2,
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(1),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_7: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(3),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(4),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_10: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(2),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(3),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_13: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(1),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(2),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_16: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(4),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(5),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_19: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(7),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(8),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_N_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_22: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(6),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(7),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_I_25: add1 port map (
      a => NN_2,
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(5),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT(6),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_IF_1_DWACT_BL_ADSBGRP0_FCI(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_1_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_iv_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_CM8I(0),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN10_AREGSIGN_SEL_M,
      S11 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_1(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_iv_1_0x: AND3A port map (
      A => GRLFPC2_0_FPI_LDOP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_1_TZ(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_iv_1_tz_0x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN5_TEMP,
      D2 => GRLFPC2_0_FPO_SIGN,
      D3 => GRLFPC2_0_FPO_SIGN,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(22),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_1_TZ(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_iv_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_1,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_IV_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_t_3_n_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N_CM8I(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC_1(0),
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_t_3_n_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_N_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_CM8I(0),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_0_0_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_1: AND3C port map (
      A => GRLFPC2_0_FPI_LDOP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(22),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN5_TEMP,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_1_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      Y => NN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_2_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_3_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_4_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_5_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_5(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_6_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_6(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_7_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_7(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_8_0x: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_0_0(0),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_8(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un4_temp_2_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      S00 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      S01 => NN_4,
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3668);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un4_temp_u_0x: CM8 port map (
      D0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(19),
      D1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3668,
      D2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN4_TEMP_U_CM8I(0),
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3668,
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5),
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
      S10 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      S11 => NN_2,
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3671);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un4_temp_u_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN4_TEMP_U_CM8I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_4: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(0),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN(0),
      s => GRLFPC2_0_FPO_EXP(0),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_7: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(9),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(9),
      s => GRLFPC2_0_FPO_EXP(9),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_10: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(5),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(5),
      s => GRLFPC2_0_FPO_EXP(5),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_13: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(1),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(1),
      s => GRLFPC2_0_FPO_EXP(1),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_16: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(10),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(10),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(10),
      s => GRLFPC2_0_FPO_EXP(10),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_19: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(6),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(6),
      s => GRLFPC2_0_FPO_EXP(6),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_22: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(2),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(2),
      s => GRLFPC2_0_FPO_EXP(2),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_25: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(11),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(11),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(11),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(11),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_28: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(7),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(7),
      s => GRLFPC2_0_FPO_EXP(7),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_31: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(3),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(3),
      s => GRLFPC2_0_FPO_EXP(3),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_34: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(12),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(12),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(12),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE(12),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_N_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_37: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(8),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(8),
      s => GRLFPC2_0_FPO_EXP(8),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_0_0_I_40: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN40_EXPXBUS(4),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(4),
      s => GRLFPC2_0_FPO_EXP(4),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_4: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(43),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(43),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(43),
      s => GRLFPC2_0_FPO_FRAC(43),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_7: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(27),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(27),
      s => GRLFPC2_0_FPO_FRAC(27),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_10: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(14),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(14),
      s => GRLFPC2_0_FPO_FRAC(14),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_13: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(1),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(1),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(1),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_16: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(28),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(28),
      s => GRLFPC2_0_FPO_FRAC(28),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_19: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(15),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(15),
      s => GRLFPC2_0_FPO_FRAC(15),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_22: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(2),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(2),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(2),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_25: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(29),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(29),
      s => GRLFPC2_0_FPO_FRAC(29),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_28: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(16),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(16),
      s => GRLFPC2_0_FPO_FRAC(16),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_31: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(3),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(3),
      s => GRLFPC2_0_FPO_FRAC(3),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_34: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(52),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(52),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(52),
      s => GRLFPC2_0_FPO_FRAC(52),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_37: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(57),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(57),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(57),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_N_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_37_0: BUFF port map (
      A => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(57),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_40: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(44),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(44),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(44),
      s => GRLFPC2_0_FPO_FRAC(44),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_43: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(12),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(12),
      s => GRLFPC2_0_FPO_FRAC(12),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_46: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(25),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(25),
      s => GRLFPC2_0_FPO_FRAC(25),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_49: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(24),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(24),
      s => GRLFPC2_0_FPO_FRAC(24),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_52: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(11),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(11),
      s => GRLFPC2_0_FPO_FRAC(11),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_55: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(38),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(38),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(38),
      s => GRLFPC2_0_FPO_FRAC(38),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_58: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(6),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(6),
      s => GRLFPC2_0_FPO_FRAC(6),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_61: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(33),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(33),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(33),
      s => GRLFPC2_0_FPO_FRAC(33),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_64: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(20),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(20),
      s => GRLFPC2_0_FPO_FRAC(20),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_67: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(7),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(7),
      s => GRLFPC2_0_FPO_FRAC(7),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_70: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(34),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(34),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(34),
      s => GRLFPC2_0_FPO_FRAC(34),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_73: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(21),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(21),
      s => GRLFPC2_0_FPO_FRAC(21),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_76: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(8),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(8),
      s => GRLFPC2_0_FPO_FRAC(8),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_79: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(35),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(35),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(35),
      s => GRLFPC2_0_FPO_FRAC(35),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_82: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(22),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(22),
      s => GRLFPC2_0_FPO_FRAC(22),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_85: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(9),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(9),
      s => GRLFPC2_0_FPO_FRAC(9),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_88: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(36),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(36),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(36),
      s => GRLFPC2_0_FPO_FRAC(36),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_91: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(23),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(23),
      s => GRLFPC2_0_FPO_FRAC(23),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_94: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(10),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(10),
      s => GRLFPC2_0_FPO_FRAC(10),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_97: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(37),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(37),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(37),
      s => GRLFPC2_0_FPO_FRAC(37),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_100: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(45),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(45),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(45),
      s => GRLFPC2_0_FPO_FRAC(45),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_103: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(48),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(48),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(48),
      s => GRLFPC2_0_FPO_FRAC(48),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_106: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(47),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(47),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(47),
      s => GRLFPC2_0_FPO_FRAC(47),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_109: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(46),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(46),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(46),
      s => GRLFPC2_0_FPO_FRAC(46),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_112: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(53),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(53),
      s => GRLFPC2_0_FPO_FRAC(53),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_115: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(30),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(30),
      s => GRLFPC2_0_FPO_FRAC(30),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_118: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(17),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(17),
      s => GRLFPC2_0_FPO_FRAC(17),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_121: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(4),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(4),
      s => GRLFPC2_0_FPO_FRAC(4),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_124: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(40),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(40),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(40),
      s => GRLFPC2_0_FPO_FRAC(40),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_127: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(49),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(49),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(49),
      s => GRLFPC2_0_FPO_FRAC(49),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_130: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(54),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(54),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(54),
      s => GRLFPC2_0_FPO_FRAC(54),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_130_0: BUFF port map (
      A => GRLFPC2_0_FPO_FRAC(54),
      Y => GRLFPC2_0_FPO_FRAC_0(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_133: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(41),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(41),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(41),
      s => GRLFPC2_0_FPO_FRAC(41),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_136: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(50),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(50),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(50),
      s => GRLFPC2_0_FPO_FRAC(50),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_139: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(55),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(55),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(55),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_142: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(42),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(42),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(42),
      s => GRLFPC2_0_FPO_FRAC(42),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_145: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(51),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(51),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(51),
      s => GRLFPC2_0_FPO_FRAC(51),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_148: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(56),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(56),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(56),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(56),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_151: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(31),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(31),
      s => GRLFPC2_0_FPO_FRAC(31),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_154: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(39),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(39),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(39),
      s => GRLFPC2_0_FPO_FRAC(39),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_157: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(26),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(26),
      s => GRLFPC2_0_FPO_FRAC(26),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_160: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(13),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(13),
      s => GRLFPC2_0_FPO_FRAC(13),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_163: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(0),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_3671,
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
      s => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF(0),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_166: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(18),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(18),
      s => GRLFPC2_0_FPO_FRAC(18),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_169: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(5),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(5),
      s => GRLFPC2_0_FPO_FRAC(5),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_172: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(32),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(32),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(32),
      s => GRLFPC2_0_FPO_FRAC(32),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf_0_0_I_175: add1 port map (
      a => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
      b => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN19_XZXBUS(19),
      fci => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(19),
      s => GRLFPC2_0_FPO_FRAC(19),
      fco => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_0_0_IF_1_DWACT_BL_ADSBGRP0_FCI(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_wqsctrl_1_68x: AND3B port map (
      A => GRLFPC2_0_FPI_LDOP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(12),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_wqsctrl_1_0_68x: AND3B port map (
      A => GRLFPC2_0_FPI_LDOP,
      B => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(12),
      C => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
      Y => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_0(68));
  x_grlfpc2_0_m7_0: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_COMB_FPDECODE_MOV2,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_M7_0_CM8I,
      S01 => cpi_d_inst(23),
      S10 => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0,
      S11 => GRLFPC2_0_COMB_FPDECODE_MOV6,
      Y => GRLFPC2_0_M7_0);
  x_grlfpc2_0_m7_0_cm8i: CM8INV port map (
      A => cpi_d_inst(19),
      Y => GRLFPC2_0_M7_0_CM8I);
  x_grlfpc2_0_m7_1: AND2A port map (
      A => cpi_d_inst(20),
      B => cpi_d_inst(21),
      Y => GRLFPC2_0_N_16_1);
  x_grlfpc2_0_m10: AND3A port map (
      A => GRLFPC2_0_COMB_FPDECODE_AFQ3_1,
      B => GRLFPC2_0_N_17_1,
      C => cpi_d_inst(20),
      Y => GRLFPC2_0_N_17);
  x_grlfpc2_0_m10_1: AND2A port map (
      A => cpi_d_inst(23),
      B => cpi_d_inst(19),
      Y => GRLFPC2_0_N_17_1);
  x_grlfpc2_0_m11: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_N_17,
      D2 => GRLFPC2_0_N_16_1,
      D3 => GRLFPC2_0_N_17,
      S00 => cpi_d_inst(30),
      S01 => NN_4,
      S10 => GRLFPC2_0_M7_0,
      S11 => NN_2,
      Y => GRLFPC2_0_N_12);
  x_grlfpc2_0_m14: AND3 port map (
      A => cpi_d_inst(31),
      B => GRLFPC2_0_COMB_RDD_1_1,
      C => GRLFPC2_0_N_12,
      Y => GRLFPC2_0_COMB_RDD_1);
  x_grlfpc2_0_m14_1: AND2A port map (
      A => cpi_d_inst(22),
      B => cpi_d_inst(24),
      Y => GRLFPC2_0_COMB_RDD_1_1);
  x_grlfpc2_0_mov_5_sqmuxa: AND3 port map (
      A => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      B => GRLFPC2_0_COMB_FPDECODE_MOV11,
      C => GRLFPC2_0_COMB_FPDECODE_MOV7,
      Y => GRLFPC2_0_MOV_5_SQMUXA);
  x_grlfpc2_0_mov_7_sqmuxa: AND2 port map (
      A => GRLFPC2_0_COMB_FPDECODE_MOV12,
      B => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      Y => GRLFPC2_0_MOV_7_SQMUXA);
  x_grlfpc2_0_op1_32x: CM8 port map (
      D0 => rfo1_data1(0),
      D1 => rfo2_data1(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(32));
  x_grlfpc2_0_op1_33x: CM8 port map (
      D0 => rfo1_data1(1),
      D1 => rfo2_data1(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(33));
  x_grlfpc2_0_op1_34x: CM8 port map (
      D0 => rfo1_data1(2),
      D1 => rfo2_data1(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(34));
  x_grlfpc2_0_op1_35x: CM8 port map (
      D0 => rfo1_data1(3),
      D1 => rfo2_data1(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(35));
  x_grlfpc2_0_op1_36x: CM8 port map (
      D0 => rfo1_data1(4),
      D1 => rfo2_data1(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(36));
  x_grlfpc2_0_op1_37x: CM8 port map (
      D0 => rfo1_data1(5),
      D1 => rfo2_data1(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(37));
  x_grlfpc2_0_op1_38x: CM8 port map (
      D0 => rfo1_data1(6),
      D1 => rfo2_data1(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(38));
  x_grlfpc2_0_op1_39x: CM8 port map (
      D0 => rfo1_data1(7),
      D1 => rfo2_data1(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(39));
  x_grlfpc2_0_op1_40x: CM8 port map (
      D0 => rfo1_data1(8),
      D1 => rfo2_data1(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(40));
  x_grlfpc2_0_op1_41x: CM8 port map (
      D0 => rfo1_data1(9),
      D1 => rfo2_data1(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(41));
  x_grlfpc2_0_op1_42x: CM8 port map (
      D0 => rfo1_data1(10),
      D1 => rfo2_data1(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(42));
  x_grlfpc2_0_op1_43x: CM8 port map (
      D0 => rfo1_data1(11),
      D1 => rfo2_data1(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(43));
  x_grlfpc2_0_op1_44x: CM8 port map (
      D0 => rfo1_data1(12),
      D1 => rfo2_data1(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(44));
  x_grlfpc2_0_op1_45x: CM8 port map (
      D0 => rfo1_data1(13),
      D1 => rfo2_data1(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(45));
  x_grlfpc2_0_op1_46x: CM8 port map (
      D0 => rfo1_data1(14),
      D1 => rfo2_data1(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(46));
  x_grlfpc2_0_op1_47x: CM8 port map (
      D0 => rfo1_data1(15),
      D1 => rfo2_data1(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(47));
  x_grlfpc2_0_op1_48x: CM8 port map (
      D0 => rfo1_data1(16),
      D1 => rfo2_data1(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(48));
  x_grlfpc2_0_op1_49x: CM8 port map (
      D0 => rfo1_data1(17),
      D1 => rfo2_data1(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(49));
  x_grlfpc2_0_op1_50x: CM8 port map (
      D0 => rfo1_data1(18),
      D1 => rfo2_data1(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(50));
  x_grlfpc2_0_op1_51x: CM8 port map (
      D0 => rfo1_data1(19),
      D1 => rfo2_data1(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(51));
  x_grlfpc2_0_op1_52x: CM8 port map (
      D0 => rfo1_data1(20),
      D1 => rfo2_data1(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(52));
  x_grlfpc2_0_op1_53x: CM8 port map (
      D0 => rfo1_data1(21),
      D1 => rfo2_data1(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(53));
  x_grlfpc2_0_op1_54x: CM8 port map (
      D0 => rfo1_data1(22),
      D1 => rfo2_data1(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(54));
  x_grlfpc2_0_op1_55x: CM8 port map (
      D0 => rfo1_data1(23),
      D1 => rfo2_data1(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(55));
  x_grlfpc2_0_op1_56x: CM8 port map (
      D0 => rfo1_data1(24),
      D1 => rfo2_data1(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(56));
  x_grlfpc2_0_op1_57x: CM8 port map (
      D0 => rfo1_data1(25),
      D1 => rfo2_data1(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(57));
  x_grlfpc2_0_op1_58x: CM8 port map (
      D0 => rfo1_data1(26),
      D1 => rfo2_data1(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(58));
  x_grlfpc2_0_op1_59x: CM8 port map (
      D0 => rfo1_data1(27),
      D1 => rfo2_data1(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(59));
  x_grlfpc2_0_op1_60x: CM8 port map (
      D0 => rfo1_data1(28),
      D1 => rfo2_data1(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(60));
  x_grlfpc2_0_op1_61x: CM8 port map (
      D0 => rfo1_data1(29),
      D1 => rfo2_data1(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(61));
  x_grlfpc2_0_op1_62x: CM8 port map (
      D0 => rfo1_data1(30),
      D1 => rfo2_data1(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(62));
  x_grlfpc2_0_op1_63x: CM8 port map (
      D0 => rfo1_data1(31),
      D1 => rfo2_data1(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_R_A_RS1_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP1(63));
  x_grlfpc2_0_op2_32x: CM8 port map (
      D0 => rfo1_data2(0),
      D1 => rfo2_data2(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(32));
  x_grlfpc2_0_op2_33x: CM8 port map (
      D0 => rfo1_data2(1),
      D1 => rfo2_data2(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(33));
  x_grlfpc2_0_op2_34x: CM8 port map (
      D0 => rfo1_data2(2),
      D1 => rfo2_data2(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(34));
  x_grlfpc2_0_op2_35x: CM8 port map (
      D0 => rfo1_data2(3),
      D1 => rfo2_data2(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(35));
  x_grlfpc2_0_op2_36x: CM8 port map (
      D0 => rfo1_data2(4),
      D1 => rfo2_data2(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(36));
  x_grlfpc2_0_op2_37x: CM8 port map (
      D0 => rfo1_data2(5),
      D1 => rfo2_data2(5),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(37));
  x_grlfpc2_0_op2_38x: CM8 port map (
      D0 => rfo1_data2(6),
      D1 => rfo2_data2(6),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(38));
  x_grlfpc2_0_op2_39x: CM8 port map (
      D0 => rfo1_data2(7),
      D1 => rfo2_data2(7),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(39));
  x_grlfpc2_0_op2_40x: CM8 port map (
      D0 => rfo1_data2(8),
      D1 => rfo2_data2(8),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(40));
  x_grlfpc2_0_op2_41x: CM8 port map (
      D0 => rfo1_data2(9),
      D1 => rfo2_data2(9),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(41));
  x_grlfpc2_0_op2_42x: CM8 port map (
      D0 => rfo1_data2(10),
      D1 => rfo2_data2(10),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(42));
  x_grlfpc2_0_op2_43x: CM8 port map (
      D0 => rfo1_data2(11),
      D1 => rfo2_data2(11),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(43));
  x_grlfpc2_0_op2_44x: CM8 port map (
      D0 => rfo1_data2(12),
      D1 => rfo2_data2(12),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(44));
  x_grlfpc2_0_op2_45x: CM8 port map (
      D0 => rfo1_data2(13),
      D1 => rfo2_data2(13),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(45));
  x_grlfpc2_0_op2_46x: CM8 port map (
      D0 => rfo1_data2(14),
      D1 => rfo2_data2(14),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(46));
  x_grlfpc2_0_op2_47x: CM8 port map (
      D0 => rfo1_data2(15),
      D1 => rfo2_data2(15),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(47));
  x_grlfpc2_0_op2_48x: CM8 port map (
      D0 => rfo1_data2(16),
      D1 => rfo2_data2(16),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(48));
  x_grlfpc2_0_op2_49x: CM8 port map (
      D0 => rfo1_data2(17),
      D1 => rfo2_data2(17),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_1,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(49));
  x_grlfpc2_0_op2_50x: CM8 port map (
      D0 => rfo1_data2(18),
      D1 => rfo2_data2(18),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(50));
  x_grlfpc2_0_op2_51x: CM8 port map (
      D0 => rfo1_data2(19),
      D1 => rfo2_data2(19),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(51));
  x_grlfpc2_0_op2_52x: CM8 port map (
      D0 => rfo1_data2(20),
      D1 => rfo2_data2(20),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(52));
  x_grlfpc2_0_op2_53x: CM8 port map (
      D0 => rfo1_data2(21),
      D1 => rfo2_data2(21),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(53));
  x_grlfpc2_0_op2_54x: CM8 port map (
      D0 => rfo1_data2(22),
      D1 => rfo2_data2(22),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(54));
  x_grlfpc2_0_op2_55x: CM8 port map (
      D0 => rfo1_data2(23),
      D1 => rfo2_data2(23),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(55));
  x_grlfpc2_0_op2_56x: CM8 port map (
      D0 => rfo1_data2(24),
      D1 => rfo2_data2(24),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(56));
  x_grlfpc2_0_op2_57x: CM8 port map (
      D0 => rfo1_data2(25),
      D1 => rfo2_data2(25),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(57));
  x_grlfpc2_0_op2_58x: CM8 port map (
      D0 => rfo1_data2(26),
      D1 => rfo2_data2(26),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4_2,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(58));
  x_grlfpc2_0_op2_59x: CM8 port map (
      D0 => rfo1_data2(27),
      D1 => rfo2_data2(27),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(59));
  x_grlfpc2_0_op2_60x: CM8 port map (
      D0 => rfo1_data2(28),
      D1 => rfo2_data2(28),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(60));
  x_grlfpc2_0_op2_61x: CM8 port map (
      D0 => rfo1_data2(29),
      D1 => rfo2_data2(29),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(61));
  x_grlfpc2_0_op2_62x: CM8 port map (
      D0 => rfo1_data2(30),
      D1 => rfo2_data2(30),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(62));
  x_grlfpc2_0_op2_63x: CM8 port map (
      D0 => rfo1_data2(31),
      D1 => rfo2_data2(31),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_UN1_FPCI_4,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_OP2(63));
  x_grlfpc2_0_r_a_afq: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFQ_1,
      E => HOLDN_I_1,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFQ);
  x_grlfpc2_0_r_a_afq_0: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFQ_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFQ_0);
  x_grlfpc2_0_r_a_afq_1: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFQ_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFQ_1);
  x_grlfpc2_0_r_a_afq_2: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFQ_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFQ_2);
  x_grlfpc2_0_r_a_afsr: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFSR_1,
      E => HOLDN_I_1,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFSR);
  x_grlfpc2_0_r_a_afsr_0: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFSR_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFSR_0);
  x_grlfpc2_0_r_a_afsr_1: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFSR_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFSR_1);
  x_grlfpc2_0_r_a_afsr_2: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_AFSR_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_AFSR_2);
  x_grlfpc2_0_r_a_fpop: DFE1B port map (
      D => GRLFPC2_0_COMB_FPOP_1,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_FPOP);
  x_grlfpc2_0_r_a_fpop_0: DFE1B port map (
      D => GRLFPC2_0_COMB_FPOP_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_A_FPOP_0);
  x_grlfpc2_0_r_a_ld: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_LD_1,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_LD);
  x_grlfpc2_0_r_a_mov: DFE1B port map (
      D => GRLFPC2_0_MOV_5_SQMUXA,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_MOV);
  x_grlfpc2_0_r_a_rdd: DFE1B port map (
      D => GRLFPC2_0_COMB_RDD_1,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RDD);
  x_grlfpc2_0_r_a_rf1ren_1x: DFE1B port map (
      D => GRLFPC2_0_N_1132,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RF1REN(1));
  x_grlfpc2_0_r_a_rf1ren_2x: DFE1B port map (
      D => GRLFPC2_0_N_1093,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RF1REN(2));
  x_grlfpc2_0_r_a_rf2ren_1x: DFE1B port map (
      D => GRLFPC2_0_N_1104,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RF2REN(1));
  x_grlfpc2_0_r_a_rf2ren_2x: DFE1B port map (
      D => GRLFPC2_0_N_1123,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RF2REN(2));
  x_grlfpc2_0_r_a_rs1_0x: DF1 port map (
      D => GRLFPC2_0_COMB_RS1_1(0),
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS1(0));
  x_grlfpc2_0_r_a_rs1_1x: DF1 port map (
      D => GRLFPC2_0_COMB_RS1_1(1),
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS1(1));
  x_grlfpc2_0_r_a_rs1_2x: DF1 port map (
      D => GRLFPC2_0_COMB_RS1_1(2),
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS1(2));
  x_grlfpc2_0_r_a_rs1_3x: DF1 port map (
      D => GRLFPC2_0_COMB_RS1_1(3),
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS1(3));
  x_grlfpc2_0_r_a_rs1_4x: DF1 port map (
      D => GRLFPC2_0_COMB_RS1_1(4),
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS1(4));
  x_grlfpc2_0_r_a_rs1d: DFE1B port map (
      D => GRLFPC2_0_COMB_RS1D_1,
      E => HOLDN_I_2,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS1D);
  x_grlfpc2_0_r_a_rs2_0x: DF1 port map (
      D => GRLFPC2_0_COMB_RS2_1(0),
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS2(0));
  x_grlfpc2_0_r_a_rs2_1x: DF1 port map (
      D => RFI2_RD2ADDR_0_INT_9_INT_22,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS2(1));
  x_grlfpc2_0_r_a_rs2_2x: DF1 port map (
      D => RFI2_RD2ADDR_1_INT_10_INT_23,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS2(2));
  x_grlfpc2_0_r_a_rs2_3x: DF1 port map (
      D => RFI2_RD2ADDR_2_INT_11_INT_24,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS2(3));
  x_grlfpc2_0_r_a_rs2_4x: DF1 port map (
      D => RFI2_RD2ADDR_3_INT_12_INT_25,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS2(4));
  x_grlfpc2_0_r_a_rs2d: DFE1B port map (
      D => GRLFPC2_0_COMB_RS2D_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_A_RS2D);
  x_grlfpc2_0_r_a_seqerr: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_SEQERR_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_A_SEQERR);
  x_grlfpc2_0_r_a_st: DFE1B port map (
      D => GRLFPC2_0_COMB_V_A_ST_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_A_ST);
  x_grlfpc2_0_r_e_afq: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_AFQ_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_E_AFQ);
  x_grlfpc2_0_r_e_afsr: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_AFSR_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_E_AFSR);
  x_grlfpc2_0_r_e_fpop: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_FPOP_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_E_FPOP);
  x_grlfpc2_0_r_e_ld: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_LD_1,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_E_LD);
  x_grlfpc2_0_r_e_rdd: DFE1B port map (
      D => GRLFPC2_0_R_A_RDD,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_E_RDD);
  x_grlfpc2_0_r_e_seqerr: DFE1B port map (
      D => GRLFPC2_0_R_A_SEQERR,
      E => HOLDN_I_3,
      CLK => clk,
      Q => GRLFPC2_0_R_E_SEQERR);
  x_grlfpc2_0_r_e_stdata_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(0),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(0));
  x_grlfpc2_0_r_e_stdata_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(1),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(1));
  x_grlfpc2_0_r_e_stdata_2x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(2),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(2));
  x_grlfpc2_0_r_e_stdata_3x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(3),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(3));
  x_grlfpc2_0_r_e_stdata_4x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(4),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(4));
  x_grlfpc2_0_r_e_stdata_5x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(5),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(5));
  x_grlfpc2_0_r_e_stdata_6x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(6),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(6));
  x_grlfpc2_0_r_e_stdata_7x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(7),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(7));
  x_grlfpc2_0_r_e_stdata_8x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(8),
      E => HOLDN_I_4,
      CLK => clk,
      Q => cpo_data(8));
  x_grlfpc2_0_r_e_stdata_9x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(9),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(9));
  x_grlfpc2_0_r_e_stdata_10x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(10),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(10));
  x_grlfpc2_0_r_e_stdata_11x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(11),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(11));
  x_grlfpc2_0_r_e_stdata_12x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(12),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(12));
  x_grlfpc2_0_r_e_stdata_13x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(13),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(13));
  x_grlfpc2_0_r_e_stdata_14x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(14),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(14));
  x_grlfpc2_0_r_e_stdata_15x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(15),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(15));
  x_grlfpc2_0_r_e_stdata_16x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(16),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(16));
  x_grlfpc2_0_r_e_stdata_17x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(17),
      E => HOLDN_I_5,
      CLK => clk,
      Q => cpo_data(17));
  x_grlfpc2_0_r_e_stdata_18x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(18),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(18));
  x_grlfpc2_0_r_e_stdata_19x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(19),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(19));
  x_grlfpc2_0_r_e_stdata_20x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(20),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(20));
  x_grlfpc2_0_r_e_stdata_21x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(21),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(21));
  x_grlfpc2_0_r_e_stdata_22x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(22),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(22));
  x_grlfpc2_0_r_e_stdata_23x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(23),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(23));
  x_grlfpc2_0_r_e_stdata_24x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(24),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(24));
  x_grlfpc2_0_r_e_stdata_25x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(25),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(25));
  x_grlfpc2_0_r_e_stdata_26x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(26),
      E => HOLDN_I_6,
      CLK => clk,
      Q => cpo_data(26));
  x_grlfpc2_0_r_e_stdata_27x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(27),
      E => HOLDN_I_7,
      CLK => clk,
      Q => cpo_data(27));
  x_grlfpc2_0_r_e_stdata_28x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(28),
      E => HOLDN_I_7,
      CLK => clk,
      Q => cpo_data(28));
  x_grlfpc2_0_r_e_stdata_29x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(29),
      E => HOLDN_I_7,
      CLK => clk,
      Q => cpo_data(29));
  x_grlfpc2_0_r_e_stdata_30x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(30),
      E => HOLDN_I_7,
      CLK => clk,
      Q => cpo_data(30));
  x_grlfpc2_0_r_e_stdata_31x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_E_STDATA_1(31),
      E => HOLDN_I_7,
      CLK => clk,
      Q => cpo_data(31));
  x_grlfpc2_0_r_fsr_aexc_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_AEXC_1(0),
      E => HOLDN_I_7,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_AEXC(0));
  x_grlfpc2_0_r_fsr_aexc_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_AEXC_1(1),
      E => HOLDN_I_7,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_AEXC(1));
  x_grlfpc2_0_r_fsr_aexc_2x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_AEXC_1(2),
      E => HOLDN_I_7,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_AEXC(2));
  x_grlfpc2_0_r_fsr_aexc_3x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_AEXC_1(3),
      E => HOLDN_I_7,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_AEXC(3));
  x_grlfpc2_0_r_fsr_aexc_4x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_AEXC_1(4),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_AEXC(4));
  x_grlfpc2_0_r_fsr_cexc_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_CEXC_1(0),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_CEXC(0));
  x_grlfpc2_0_r_fsr_cexc_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_CEXC_1(1),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_CEXC(1));
  x_grlfpc2_0_r_fsr_cexc_2x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_CEXC_1(2),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_CEXC(2));
  x_grlfpc2_0_r_fsr_cexc_3x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_CEXC_1(3),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_CEXC(3));
  x_grlfpc2_0_r_fsr_cexc_4x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_CEXC_1(4),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_CEXC(4));
  x_grlfpc2_0_r_fsr_fcc_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_FCC_1(0),
      E => HOLDN_I_8,
      CLK => clk,
      Q => CPO_CC_0_INT_2);
  x_grlfpc2_0_r_fsr_fcc_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_FCC_1(1),
      E => HOLDN_I_8,
      CLK => clk,
      Q => CPO_CC_1_INT_3);
  x_grlfpc2_0_r_fsr_ftt_0x: DFE1B port map (
      D => GRLFPC2_0_V_FSR_FTT_1(0),
      E => HOLDN_I_8,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_FTT(0));
  x_grlfpc2_0_r_fsr_ftt_2x: DFE1B port map (
      D => GRLFPC2_0_V_FSR_FTT_1(2),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_FTT(2));
  x_grlfpc2_0_r_fsr_nonstd: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_NONSTD_1,
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_NONSTD);
  x_grlfpc2_0_r_fsr_rd_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_RD_1(0),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_RD(0));
  x_grlfpc2_0_r_fsr_rd_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_RD_1(1),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_RD(1));
  x_grlfpc2_0_r_fsr_tem_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(0),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_TEM(0));
  x_grlfpc2_0_r_fsr_tem_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(1),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_TEM(1));
  x_grlfpc2_0_r_fsr_tem_2x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(2),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_TEM(2));
  x_grlfpc2_0_r_fsr_tem_3x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(3),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_TEM(3));
  x_grlfpc2_0_r_fsr_tem_4x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(4),
      E => HOLDN_I_9,
      CLK => clk,
      Q => GRLFPC2_0_R_FSR_TEM(4));
  x_grlfpc2_0_r_i_cc_0x: DFE1B port map (
      D => GRLFPC2_0_FPO_CC(0),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      CLK => clk,
      Q => GRLFPC2_0_R_I_CC(0));
  x_grlfpc2_0_r_i_cc_1x: DFE1B port map (
      D => GRLFPC2_0_FPO_CC(1),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      CLK => clk,
      Q => GRLFPC2_0_R_I_CC(1));
  x_grlfpc2_0_r_i_exc_0x: DF1 port map (
      D => GRLFPC2_0_N_163,
      CLK => clk,
      Q => GRLFPC2_0_R_I_EXC(0));
  x_grlfpc2_0_r_i_exc_1x: DF1 port map (
      D => GRLFPC2_0_N_164,
      CLK => clk,
      Q => GRLFPC2_0_R_I_EXC(1));
  x_grlfpc2_0_r_i_exc_2x: DF1 port map (
      D => GRLFPC2_0_N_165,
      CLK => clk,
      Q => GRLFPC2_0_R_I_EXC(2));
  x_grlfpc2_0_r_i_exc_3x: DF1 port map (
      D => GRLFPC2_0_N_166,
      CLK => clk,
      Q => GRLFPC2_0_R_I_EXC(3));
  x_grlfpc2_0_r_i_exc_4x: DF1 port map (
      D => GRLFPC2_0_N_167,
      CLK => clk,
      Q => GRLFPC2_0_R_I_EXC(4));
  x_grlfpc2_0_r_i_exc_1_0x: CM8 port map (
      D0 => GRLFPC2_0_R_I_EXC(0),
      D1 => GRLFPC2_0_FPO_EXC(0),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_UN1_HOLDN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN_3,
      S11 => NN_2,
      Y => GRLFPC2_0_N_163);
  x_grlfpc2_0_r_i_exc_1_1x: CM8 port map (
      D0 => GRLFPC2_0_R_I_EXC(1),
      D1 => GRLFPC2_0_FPO_EXC(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_UN1_HOLDN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN,
      S11 => NN_2,
      Y => GRLFPC2_0_N_164);
  x_grlfpc2_0_r_i_exc_1_2x: CM8 port map (
      D0 => GRLFPC2_0_R_I_EXC(2),
      D1 => GRLFPC2_0_R_I_EXC(2),
      D2 => NN_2,
      D3 => GRLFPC2_0_FPO_EXC(0),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_0(2),
      S01 => GRLFPC2_0_R_I_EXC_1_CM8I(2),
      S10 => GRLFPC2_0_COMB_UN2_HOLDN,
      S11 => GRLFPC2_0_UN1_HOLDN_1,
      Y => GRLFPC2_0_N_165);
  x_grlfpc2_0_r_i_exc_1_3x: CM8 port map (
      D0 => GRLFPC2_0_R_I_EXC(3),
      D1 => GRLFPC2_0_FPO_EXC(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_UN1_HOLDN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN,
      S11 => NN_2,
      Y => GRLFPC2_0_N_166);
  x_grlfpc2_0_r_i_exc_1_4x: CM8 port map (
      D0 => GRLFPC2_0_R_I_EXC(4),
      D1 => GRLFPC2_0_FPO_EXC(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_UN1_HOLDN_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_COMB_UN2_HOLDN,
      S11 => NN_2,
      Y => GRLFPC2_0_N_167);
  x_grlfpc2_0_r_i_exc_1_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_COMB_UN2_HOLDN,
      Y => GRLFPC2_0_R_I_EXC_1_CM8I(2));
  x_grlfpc2_0_r_i_exec: DFE1B port map (
      D => GRLFPC2_0_N_1063,
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_EXEC);
  x_grlfpc2_0_r_i_inst_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(0),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(0));
  x_grlfpc2_0_r_i_inst_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(1),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(1));
  x_grlfpc2_0_r_i_inst_2x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(2),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(2));
  x_grlfpc2_0_r_i_inst_3x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(3),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(3));
  x_grlfpc2_0_r_i_inst_4x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(4),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(4));
  x_grlfpc2_0_r_i_inst_5x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(5),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(5));
  x_grlfpc2_0_r_i_inst_6x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(6),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(6));
  x_grlfpc2_0_r_i_inst_7x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(7),
      E => HOLDN_I_10,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(7));
  x_grlfpc2_0_r_i_inst_8x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(8),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(8));
  x_grlfpc2_0_r_i_inst_9x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(9),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(9));
  x_grlfpc2_0_r_i_inst_10x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(10),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(10));
  x_grlfpc2_0_r_i_inst_11x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(11),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(11));
  x_grlfpc2_0_r_i_inst_12x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(12),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(12));
  x_grlfpc2_0_r_i_inst_13x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(13),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(13));
  x_grlfpc2_0_r_i_inst_14x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(14),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(14));
  x_grlfpc2_0_r_i_inst_15x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(15),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(15));
  x_grlfpc2_0_r_i_inst_16x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(16),
      E => HOLDN_I_11,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(16));
  x_grlfpc2_0_r_i_inst_17x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(17),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(17));
  x_grlfpc2_0_r_i_inst_18x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(18),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(18));
  x_grlfpc2_0_r_i_inst_19x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(19),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(19));
  x_grlfpc2_0_r_i_inst_20x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(20),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(20));
  x_grlfpc2_0_r_i_inst_21x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(21),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(21));
  x_grlfpc2_0_r_i_inst_22x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(22),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(22));
  x_grlfpc2_0_r_i_inst_23x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(23),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(23));
  x_grlfpc2_0_r_i_inst_24x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(24),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(24));
  x_grlfpc2_0_r_i_inst_25x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(25),
      E => HOLDN_I_12,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(25));
  x_grlfpc2_0_r_i_inst_26x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(26),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(26));
  x_grlfpc2_0_r_i_inst_27x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(27),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(27));
  x_grlfpc2_0_r_i_inst_28x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(28),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(28));
  x_grlfpc2_0_r_i_inst_29x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(29),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(29));
  x_grlfpc2_0_r_i_inst_30x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(30),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(30));
  x_grlfpc2_0_r_i_inst_31x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_INST_1(31),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_INST(31));
  x_grlfpc2_0_r_i_pc_2x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(2),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(2));
  x_grlfpc2_0_r_i_pc_3x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(3),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(3));
  x_grlfpc2_0_r_i_pc_4x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(4),
      E => HOLDN_I_13,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(4));
  x_grlfpc2_0_r_i_pc_5x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(5),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(5));
  x_grlfpc2_0_r_i_pc_6x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(6),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(6));
  x_grlfpc2_0_r_i_pc_7x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(7),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(7));
  x_grlfpc2_0_r_i_pc_8x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(8),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(8));
  x_grlfpc2_0_r_i_pc_9x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(9),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(9));
  x_grlfpc2_0_r_i_pc_10x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(10),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(10));
  x_grlfpc2_0_r_i_pc_11x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(11),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(11));
  x_grlfpc2_0_r_i_pc_12x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(12),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(12));
  x_grlfpc2_0_r_i_pc_13x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(13),
      E => HOLDN_I_14,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(13));
  x_grlfpc2_0_r_i_pc_14x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(14),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(14));
  x_grlfpc2_0_r_i_pc_15x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(15),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(15));
  x_grlfpc2_0_r_i_pc_16x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(16),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(16));
  x_grlfpc2_0_r_i_pc_17x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(17),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(17));
  x_grlfpc2_0_r_i_pc_18x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(18),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(18));
  x_grlfpc2_0_r_i_pc_19x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(19),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(19));
  x_grlfpc2_0_r_i_pc_20x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(20),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(20));
  x_grlfpc2_0_r_i_pc_21x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(21),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(21));
  x_grlfpc2_0_r_i_pc_22x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(22),
      E => HOLDN_I_15,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(22));
  x_grlfpc2_0_r_i_pc_23x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(23),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(23));
  x_grlfpc2_0_r_i_pc_24x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(24),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(24));
  x_grlfpc2_0_r_i_pc_25x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(25),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(25));
  x_grlfpc2_0_r_i_pc_26x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(26),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(26));
  x_grlfpc2_0_r_i_pc_27x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(27),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(27));
  x_grlfpc2_0_r_i_pc_28x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(28),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(28));
  x_grlfpc2_0_r_i_pc_29x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(29),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(29));
  x_grlfpc2_0_r_i_pc_30x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(30),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(30));
  x_grlfpc2_0_r_i_pc_31x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_I_PC_1(31),
      E => HOLDN_I_16,
      CLK => clk,
      Q => GRLFPC2_0_R_I_PC(31));
  x_grlfpc2_0_r_i_rdd: DFE1B port map (
      D => GRLFPC2_0_N_1080,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RDD);
  x_grlfpc2_0_r_i_res_0x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(3),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(0));
  x_grlfpc2_0_r_i_res_1x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(4),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(1));
  x_grlfpc2_0_r_i_res_2x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(5),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(2));
  x_grlfpc2_0_r_i_res_3x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(6),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(3));
  x_grlfpc2_0_r_i_res_4x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(7),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(4));
  x_grlfpc2_0_r_i_res_5x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(8),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(5));
  x_grlfpc2_0_r_i_res_6x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(9),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(6));
  x_grlfpc2_0_r_i_res_7x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(10),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(7));
  x_grlfpc2_0_r_i_res_8x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(11),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(8));
  x_grlfpc2_0_r_i_res_9x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(12),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_1,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(9));
  x_grlfpc2_0_r_i_res_10x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(13),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(10));
  x_grlfpc2_0_r_i_res_11x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(14),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(11));
  x_grlfpc2_0_r_i_res_12x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(15),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(12));
  x_grlfpc2_0_r_i_res_13x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(16),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(13));
  x_grlfpc2_0_r_i_res_14x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(17),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(14));
  x_grlfpc2_0_r_i_res_15x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(18),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(15));
  x_grlfpc2_0_r_i_res_16x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(19),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(16));
  x_grlfpc2_0_r_i_res_17x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(20),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(17));
  x_grlfpc2_0_r_i_res_18x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(21),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_2,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(18));
  x_grlfpc2_0_r_i_res_19x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(22),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(19));
  x_grlfpc2_0_r_i_res_20x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(23),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(20));
  x_grlfpc2_0_r_i_res_21x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(24),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(21));
  x_grlfpc2_0_r_i_res_22x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(25),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(22));
  x_grlfpc2_0_r_i_res_23x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(26),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(23));
  x_grlfpc2_0_r_i_res_24x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(27),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(24));
  x_grlfpc2_0_r_i_res_25x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(28),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(25));
  x_grlfpc2_0_r_i_res_26x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(29),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(26));
  x_grlfpc2_0_r_i_res_27x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(30),
      E => GRLFPC2_0_COMB_UN6_IUEXEC_3,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(27));
  x_grlfpc2_0_r_i_res_28x: DFE1B port map (
      D => GRLFPC2_0_FPO_FRAC(31),
      E => GRLFPC2_0_COMB_UN6_IUEXEC,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(28));
  x_grlfpc2_0_r_i_res_29x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(29),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(29));
  x_grlfpc2_0_r_i_res_30x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(30),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(30));
  x_grlfpc2_0_r_i_res_31x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(31),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(31));
  x_grlfpc2_0_r_i_res_32x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(32),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(32));
  x_grlfpc2_0_r_i_res_33x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(33),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(33));
  x_grlfpc2_0_r_i_res_34x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(34),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(34));
  x_grlfpc2_0_r_i_res_35x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(35),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(35));
  x_grlfpc2_0_r_i_res_36x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(36),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(36));
  x_grlfpc2_0_r_i_res_37x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(37),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(37));
  x_grlfpc2_0_r_i_res_38x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(38),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(38));
  x_grlfpc2_0_r_i_res_39x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(39),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(39));
  x_grlfpc2_0_r_i_res_40x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(40),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(40));
  x_grlfpc2_0_r_i_res_41x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(41),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(41));
  x_grlfpc2_0_r_i_res_42x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(42),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(42));
  x_grlfpc2_0_r_i_res_43x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(43),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(43));
  x_grlfpc2_0_r_i_res_44x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(44),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(44));
  x_grlfpc2_0_r_i_res_45x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(45),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(45));
  x_grlfpc2_0_r_i_res_46x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(46),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(46));
  x_grlfpc2_0_r_i_res_47x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(47),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(47));
  x_grlfpc2_0_r_i_res_48x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(48),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(48));
  x_grlfpc2_0_r_i_res_49x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(49),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(49));
  x_grlfpc2_0_r_i_res_50x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(50),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(50));
  x_grlfpc2_0_r_i_res_51x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(51),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(51));
  x_grlfpc2_0_r_i_res_52x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(52),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(52));
  x_grlfpc2_0_r_i_res_53x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(53),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(53));
  x_grlfpc2_0_r_i_res_54x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(54),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(54));
  x_grlfpc2_0_r_i_res_55x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(55),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(55));
  x_grlfpc2_0_r_i_res_56x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(56),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(56));
  x_grlfpc2_0_r_i_res_57x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(57),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(57));
  x_grlfpc2_0_r_i_res_58x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(58),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(58));
  x_grlfpc2_0_r_i_res_59x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(59),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(59));
  x_grlfpc2_0_r_i_res_60x: DFE1B port map (
      D => GRLFPC2_0_FPO_EXP(8),
      E => GRLFPC2_0_COMB_UN6_IUEXEC,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(60));
  x_grlfpc2_0_r_i_res_61x: DFE1B port map (
      D => GRLFPC2_0_FPO_EXP(9),
      E => GRLFPC2_0_COMB_UN6_IUEXEC,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(61));
  x_grlfpc2_0_r_i_res_62x: DFE1B port map (
      D => GRLFPC2_0_FPO_EXP(10),
      E => GRLFPC2_0_COMB_UN6_IUEXEC,
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(62));
  x_grlfpc2_0_r_i_res_63x: DF1 port map (
      D => GRLFPC2_0_COMB_V_I_RES_1(63),
      CLK => clk,
      Q => GRLFPC2_0_R_I_RES(63));
  x_grlfpc2_0_r_i_v: DF1 port map (
      D => GRLFPC2_0_N_169,
      CLK => clk,
      Q => GRLFPC2_0_R_I_V);
  x_grlfpc2_0_r_i_v_0: CM8 port map (
      D0 => GRLFPC2_0_COMB_V_I_V_1,
      D1 => GRLFPC2_0_R_I_V,
      D2 => GRLFPC2_0_COMB_V_I_V_1,
      D3 => GRLFPC2_0_COMB_V_I_V_1,
      S00 => GRLFPC2_0_V_I_V_1_SQMUXA,
      S01 => GRLFPC2_0_N_1063_3,
      S10 => GRLFPC2_0_COMB_V_I_V6,
      S11 => NN_2,
      Y => GRLFPC2_0_N_1);
  x_grlfpc2_0_r_i_v_1: AND2A port map (
      A => RST_I,
      B => GRLFPC2_0_N_1,
      Y => GRLFPC2_0_N_169);
  x_grlfpc2_0_r_m_afq: DFE1B port map (
      D => GRLFPC2_0_COMB_V_M_AFQ_1,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_M_AFQ);
  x_grlfpc2_0_r_m_afsr: DFE1B port map (
      D => GRLFPC2_0_COMB_V_M_AFSR_1,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_M_AFSR);
  x_grlfpc2_0_r_m_fpop: DFE1B port map (
      D => GRLFPC2_0_COMB_V_M_FPOP_1,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_M_FPOP);
  x_grlfpc2_0_r_m_ld: DFE1B port map (
      D => GRLFPC2_0_COMB_V_M_LD_1,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_M_LD);
  x_grlfpc2_0_r_m_rdd: DFE1B port map (
      D => GRLFPC2_0_R_E_RDD,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_M_RDD);
  x_grlfpc2_0_r_m_seqerr: DFE1B port map (
      D => GRLFPC2_0_R_E_SEQERR,
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_M_SEQERR);
  x_grlfpc2_0_r_mk_busy: DF1 port map (
      D => GRLFPC2_0_N_171,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_BUSY);
  x_grlfpc2_0_r_mk_busy2: DF1 port map (
      D => GRLFPC2_0_N_173,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_BUSY2);
  x_grlfpc2_0_r_mk_busy2_0: AND3B port map (
      A => GRLFPC2_0_COMB_ANNULFPU_1,
      B => RST_I,
      C => GRLFPC2_0_R_MK_BUSY,
      Y => GRLFPC2_0_N_173);
  x_grlfpc2_0_r_mk_busy_0: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => NN_4,
      D3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
      S00 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3,
      S01 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1,
      S10 => GRLFPC2_0_R_MK_BUSY_0_2,
      S11 => NN_2,
      Y => GRLFPC2_0_N_171);
  x_grlfpc2_0_r_mk_busy_0_2: AND4C port map (
      A => GRLFPC2_0_COMB_ANNULFPU_1,
      B => RST_I,
      C => GRLFPC2_0_COMB_UN10_IUEXEC,
      D => CPO_HOLDN_INT_4,
      Y => GRLFPC2_0_R_MK_BUSY_0_2);
  x_grlfpc2_0_r_mk_holdn1: DF1 port map (
      D => GRLFPC2_0_N_161,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_HOLDN1);
  x_grlfpc2_0_r_mk_holdn1_0: OR2A port map (
      A => GRLFPC2_0_R_MK_RST2,
      B => RST_I,
      Y => GRLFPC2_0_N_161);
  x_grlfpc2_0_r_mk_holdn2: DF1 port map (
      D => GRLFPC2_0_R_MK_HOLDN1,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_HOLDN2);
  x_grlfpc2_0_r_mk_ldop: DF1 port map (
      D => GRLFPC2_0_COMB_V_MK_LDOP_1,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_LDOP);
  x_grlfpc2_0_r_mk_rst: DF1 port map (
      D => GRLFPC2_0_COMB_V_MK_RST_1,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_RST);
  x_grlfpc2_0_r_mk_rst2: DF1 port map (
      D => GRLFPC2_0_R_MK_RST,
      CLK => clk,
      Q => GRLFPC2_0_R_MK_RST2);
  x_grlfpc2_0_r_state_0x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_STATE_1(0),
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_STATE(0));
  x_grlfpc2_0_r_state_1x: DFE1B port map (
      D => GRLFPC2_0_COMB_V_STATE_1(1),
      E => HOLDN_I_17,
      CLK => clk,
      Q => GRLFPC2_0_R_STATE(1));
  x_grlfpc2_0_r_x_afq: DFE1B port map (
      D => GRLFPC2_0_COMB_V_X_AFQ_1,
      E => HOLDN_I_0_1,
      CLK => clk,
      Q => GRLFPC2_0_R_X_AFQ);
  x_grlfpc2_0_r_x_afsr: DFE1B port map (
      D => GRLFPC2_0_COMB_V_X_AFSR_1,
      E => HOLDN_I,
      CLK => clk,
      Q => GRLFPC2_0_R_X_AFSR);
  x_grlfpc2_0_r_x_fpop: DFE1B port map (
      D => GRLFPC2_0_COMB_V_X_FPOP_1,
      E => HOLDN_I,
      CLK => clk,
      Q => GRLFPC2_0_R_X_FPOP);
  x_grlfpc2_0_r_x_fpop_0: DFE1B port map (
      D => GRLFPC2_0_COMB_V_X_FPOP_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_X_FPOP_0);
  x_grlfpc2_0_r_x_ld: DFE1B port map (
      D => GRLFPC2_0_COMB_V_X_LD_1,
      E => HOLDN_I,
      CLK => clk,
      Q => GRLFPC2_0_R_X_LD);
  x_grlfpc2_0_r_x_ld_0: DFE1B port map (
      D => GRLFPC2_0_COMB_V_X_LD_1,
      E => HOLDN_I_0,
      CLK => clk,
      Q => GRLFPC2_0_R_X_LD_0);
  x_grlfpc2_0_r_x_rdd: DFE1B port map (
      D => GRLFPC2_0_R_M_RDD,
      E => HOLDN_I,
      CLK => clk,
      Q => GRLFPC2_0_R_X_RDD);
  x_grlfpc2_0_r_x_seqerr: DFE1B port map (
      D => GRLFPC2_0_R_M_SEQERR,
      E => HOLDN_I,
      CLK => clk,
      Q => GRLFPC2_0_R_X_SEQERR);
  x_grlfpc2_0_rf1ren_1x: CM8 port map (
      D0 => GRLFPC2_0_N_1132_1_N,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_RF1REN_CM8I(1),
      S01 => GRLFPC2_0_COMB_RS1_1(0),
      S10 => GRLFPC2_0_R_A_RF1REN(1),
      S11 => CPI_DBG_ENABLE_0,
      Y => rfi1_ren1);
  x_grlfpc2_0_rf1ren_2x: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      D1 => NN_2,
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_RF1REN_CM8I(2),
      S01 => GRLFPC2_0_COMB_RS2_1(0),
      S10 => GRLFPC2_0_R_A_RF1REN(2),
      S11 => CPI_DBG_ENABLE_0,
      Y => rfi1_ren2);
  x_grlfpc2_0_rf1ren_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_COMB_RS1D_1,
      Y => GRLFPC2_0_RF1REN_CM8I(1));
  x_grlfpc2_0_rf1ren_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_N_1127,
      Y => GRLFPC2_0_RF1REN_CM8I(2));
  x_grlfpc2_0_rf2ren_1x: CM8 port map (
      D0 => GRLFPC2_0_N_1132_1_N,
      D1 => GRLFPC2_0_COMB_RS1_1(0),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_RF2REN_CM8I(1),
      S01 => GRLFPC2_0_N_1132_1_N,
      S10 => GRLFPC2_0_R_A_RF2REN(1),
      S11 => CPI_DBG_ENABLE_0,
      Y => rfi2_ren1);
  x_grlfpc2_0_rf2ren_2x: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      D1 => GRLFPC2_0_COMB_RS2_1(0),
      D2 => NN_4,
      D3 => NN_4,
      S00 => GRLFPC2_0_RF2REN_CM8I(2),
      S01 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      S10 => GRLFPC2_0_R_A_RF2REN(2),
      S11 => CPI_DBG_ENABLE_0,
      Y => rfi2_ren2);
  x_grlfpc2_0_rf2ren_cm8i_1x: CM8INV port map (
      A => GRLFPC2_0_COMB_RS1D_1,
      Y => GRLFPC2_0_RF2REN_CM8I(1));
  x_grlfpc2_0_rf2ren_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_N_1127,
      Y => GRLFPC2_0_RF2REN_CM8I(2));
  x_grlfpc2_0_rs1_1_1x: CM8 port map (
      D0 => GRLFPC2_0_COMB_RS1_1(1),
      D1 => cpi_dbg_addr(1),
      D2 => NN_2,
      D3 => NN_2,
      S00 => CPI_DBG_ENABLE_0,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => RFI2_RD1ADDR_0_INT_5_INT_18);
  x_grlfpc2_0_rs1_1_2x: CM8 port map (
      D0 => GRLFPC2_0_COMB_RS1_1(2),
      D1 => cpi_dbg_addr(2),
      D2 => NN_2,
      D3 => NN_2,
      S00 => cpi_dbg_enable,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => RFI2_RD1ADDR_1_INT_6_INT_19);
  x_grlfpc2_0_rs1_1_3x: CM8 port map (
      D0 => GRLFPC2_0_COMB_RS1_1(3),
      D1 => cpi_dbg_addr(3),
      D2 => NN_2,
      D3 => NN_2,
      S00 => cpi_dbg_enable,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => RFI2_RD1ADDR_2_INT_7_INT_20);
  x_grlfpc2_0_rs1_1_4x: CM8 port map (
      D0 => GRLFPC2_0_COMB_RS1_1(4),
      D1 => cpi_dbg_addr(4),
      D2 => NN_2,
      D3 => NN_2,
      S00 => cpi_dbg_enable,
      S01 => NN_4,
      S10 => NN_2,
      S11 => NN_2,
      Y => RFI2_RD1ADDR_3_INT_8_INT_21);
  x_grlfpc2_0_rs1d_cnst_0_a2: AND3 port map (
      A => cpi_d_inst(21),
      B => GRLFPC2_0_RS1D_CNST_0_A2_0,
      C => cpi_d_inst(31),
      Y => GRLFPC2_0_RS1D_CNST);
  x_grlfpc2_0_rs1d_cnst_0_a2_0: AND2 port map (
      A => GRLFPC2_0_COMB_RDD_1_1,
      B => GRLFPC2_0_N_335,
      Y => GRLFPC2_0_RS1D_CNST_0_A2_0);
  x_grlfpc2_0_rs1d_cnst_0_a3_0_0_0_n: OR2A port map (
      A => GRLFPC2_0_COMB_FPDECODE_MOV5,
      B => cpi_d_inst(30),
      Y => GRLFPC2_0_RS1D_CNST_0_A3_0_0_N);
  x_grlfpc2_0_rs1d_cnst_0_o2: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => cpi_d_inst(23),
      D3 => cpi_d_inst(30),
      S00 => cpi_d_inst(20),
      S01 => NN_4,
      S10 => GRLFPC2_0_RS1D_CNST_0_O2_CM8I,
      S11 => GRLFPC2_0_N_17_1,
      Y => GRLFPC2_0_N_335);
  x_grlfpc2_0_rs1d_cnst_0_o2_cm8i: CM8INV port map (
      A => GRLFPC2_0_RS1D_CNST_0_A3_0_0_N,
      Y => GRLFPC2_0_RS1D_CNST_0_O2_CM8I);
  x_grlfpc2_0_rs1v10: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_AFQ3,
      D1 => NN_4,
      D2 => GRLFPC2_0_COMB_FPDECODE_AFQ3,
      D3 => GRLFPC2_0_COMB_FPDECODE_AFQ3,
      S00 => GRLFPC2_0_COMB_RDD_1_1,
      S01 => GRLFPC2_0_COMB_FPDECODE_ST_1,
      S10 => cpi_d_inst(20),
      S11 => cpi_d_inst(19),
      Y => GRLFPC2_0_RS1V10);
  x_grlfpc2_0_rs1v_0_sqmuxa_1: AND2 port map (
      A => GRLFPC2_0_RS1V10,
      B => GRLFPC2_0_COMB_FPDECODE_AFQ13,
      Y => GRLFPC2_0_RS1V_0_SQMUXA_1);
  x_grlfpc2_0_rs2_0_sqmuxa: AND2 port map (
      A => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
      B => GRLFPC2_0_COMB_FPDECODE_AFQ12,
      Y => GRLFPC2_0_RS2_0_SQMUXA);
  x_grlfpc2_0_un1_fpci_2_n: CM8 port map (
      D0 => GRLFPC2_0_V_FSR_FTT_0_SQMUXA_2_1,
      D1 => GRLFPC2_0_UN1_FPCI_2_N_CM8I,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_X_AFQ,
      S01 => GRLFPC2_0_COMB_QNE2,
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_UN1_FPCI_2_N);
  x_grlfpc2_0_un1_fpci_2_n_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      Y => GRLFPC2_0_UN1_FPCI_2_N_CM8I);
  x_grlfpc2_0_un1_fpci_3_0: CM8 port map (
      D0 => GRLFPC2_0_UN1_FPCI_3_1,
      D1 => NN_4,
      D2 => GRLFPC2_0_UN1_FPCI_3_1,
      D3 => GRLFPC2_0_UN1_FPCI_3_1,
      S00 => cpi_x_inst(20),
      S01 => GRLFPC2_0_R_X_LD_0,
      S10 => GRLFPC2_0_COMB_WREN22,
      S11 => GRLFPC2_0_R_X_AFSR,
      Y => GRLFPC2_0_UN1_FPCI_3_0);
  x_grlfpc2_0_un1_fpci_3_1: OR2 port map (
      A => GRLFPC2_0_R_X_SEQERR,
      B => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      Y => GRLFPC2_0_UN1_FPCI_3_1);
  x_grlfpc2_0_un1_holdn_1: OR2A port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC,
      B => GRLFPC2_0_COMB_UN2_HOLDN,
      Y => GRLFPC2_0_UN1_HOLDN_1);
  x_grlfpc2_0_un1_holdn_1_0: OR2A port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      B => GRLFPC2_0_COMB_UN2_HOLDN_0,
      Y => GRLFPC2_0_UN1_HOLDN_1_0);
  x_grlfpc2_0_un1_holdn_1_1: OR2A port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      B => GRLFPC2_0_COMB_UN2_HOLDN_0,
      Y => GRLFPC2_0_UN1_HOLDN_1_1);
  x_grlfpc2_0_un1_holdn_1_2: OR2A port map (
      A => GRLFPC2_0_COMB_UN6_IUEXEC_0_0,
      B => GRLFPC2_0_COMB_UN2_HOLDN_0,
      Y => GRLFPC2_0_UN1_HOLDN_1_2);
  x_grlfpc2_0_un1_mov_1_sqmuxa_tz_0: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_MOV4_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_COMB_FPDECODE_MOV5,
      S01 => NN_4,
      S10 => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0_CM8I,
      S11 => cpi_d_inst(11),
      Y => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0);
  x_grlfpc2_0_un1_mov_1_sqmuxa_tz_0_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_FPDECODE_MOV4_3,
      Y => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0_CM8I);
  x_grlfpc2_0_un1_mov_1_sqmuxa_tz_1: CM8 port map (
      D0 => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_1_0,
      D1 => NN_4,
      D2 => NN_2,
      D3 => NN_4,
      S00 => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_0,
      S01 => NN_4,
      S10 => cpi_d_inst(8),
      S11 => NN_2,
      Y => GRLFPC2_0_UN1_MOV_1_SQMUXA_TZ_1);
  x_grlfpc2_0_un1_wren1_0_sqmuxa: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_WREN1_0_SQMUXA_2,
      D3 => NN_2,
      S00 => NN_2,
      S01 => NN_2,
      S10 => GRLFPC2_0_UN1_WREN1_0_SQMUXA_CM8I,
      S11 => GRLFPC2_0_UN1_FPCI_3_1,
      Y => GRLFPC2_0_UN1_WREN1_0_SQMUXA);
  x_grlfpc2_0_un1_wren1_0_sqmuxa_cm8i: CM8INV port map (
      A => GRLFPC2_0_UN1_FPCI_3_0,
      Y => GRLFPC2_0_UN1_WREN1_0_SQMUXA_CM8I);
  x_grlfpc2_0_v_fsr_ftt_0_sqmuxa_2_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      B => GRLFPC2_0_R_X_SEQERR,
      Y => GRLFPC2_0_V_FSR_FTT_0_SQMUXA_2_1);
  x_grlfpc2_0_v_fsr_ftt_1_0x: CM8 port map (
      D0 => rst,
      D1 => NN_2,
      D2 => rst,
      D3 => GRLFPC2_0_R_FSR_FTT(0),
      S00 => rst,
      S01 => GRLFPC2_0_V_FSR_FTT_1_CM8I(0),
      S10 => GRLFPC2_0_COMB_UN1_FPCI,
      S11 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA,
      Y => GRLFPC2_0_V_FSR_FTT_1(0));
  x_grlfpc2_0_v_fsr_ftt_1_2x: CM8 port map (
      D0 => NN_2,
      D1 => GRLFPC2_0_V_FSR_FTT_0_SQMUXA_2_1,
      D2 => NN_2,
      D3 => GRLFPC2_0_R_FSR_FTT(2),
      S00 => rst,
      S01 => GRLFPC2_0_V_FSR_FTT_1_CM8I(2),
      S10 => GRLFPC2_0_COMB_UN1_FPCI,
      S11 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA,
      Y => GRLFPC2_0_V_FSR_FTT_1(2));
  x_grlfpc2_0_v_fsr_ftt_1_cm8i_0x: CM8INV port map (
      A => GRLFPC2_0_COMB_V_I_V6,
      Y => GRLFPC2_0_V_FSR_FTT_1_CM8I(0));
  x_grlfpc2_0_v_fsr_ftt_1_cm8i_2x: CM8INV port map (
      A => GRLFPC2_0_COMB_V_I_V6,
      Y => GRLFPC2_0_V_FSR_FTT_1_CM8I(2));
  x_grlfpc2_0_v_fsr_ftt_1_sqmuxa: CM8 port map (
      D0 => NN_2,
      D1 => NN_4,
      D2 => NN_2,
      D3 => GRLFPC2_0_R_X_LD_0,
      S00 => GRLFPC2_0_V_STATE_1_SQMUXA_1,
      S01 => NN_4,
      S10 => GRLFPC2_0_R_X_AFSR,
      S11 => NN_2,
      Y => GRLFPC2_0_V_FSR_FTT_1_SQMUXA);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa: AND2 port map (
      A => GRLFPC2_0_R_X_LD,
      B => GRLFPC2_0_R_X_AFSR,
      Y => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_1: AND3 port map (
      A => cpi_dbg_enable,
      B => cpi_dbg_write,
      C => cpi_dbg_fsr,
      Y => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_1_0: AND3 port map (
      A => CPI_DBG_ENABLE_0,
      B => cpi_dbg_write,
      C => CPI_DBG_FSR_0,
      Y => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1_0);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_2: AND3A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI,
      B => GRLFPC2_0_R_X_LD,
      C => GRLFPC2_0_R_X_AFSR,
      Y => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_2_0: AND3A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_1_0,
      B => GRLFPC2_0_R_X_LD_0,
      C => GRLFPC2_0_R_X_AFSR,
      Y => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_0);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_2_1: AND3A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_LD_0,
      C => GRLFPC2_0_R_X_AFSR,
      Y => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_2_1);
  x_grlfpc2_0_v_i_exec_0_sqmuxa: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI,
      B => GRLFPC2_0_R_X_FPOP,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_0: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_0);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_1: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_1);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_2: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_2);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_3: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_3);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_4: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_4);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_5: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_5);
  x_grlfpc2_0_v_i_exec_0_sqmuxa_6: AND2A port map (
      A => GRLFPC2_0_COMB_UN1_FPCI_0,
      B => GRLFPC2_0_R_X_FPOP_0,
      Y => GRLFPC2_0_V_I_EXEC_0_SQMUXA_6);
  x_grlfpc2_0_v_i_v_1_sqmuxa: AND3B port map (
      A => GRLFPC2_0_COMB_ANNULRES_1,
      B => GRLFPC2_0_COMB_UN2_HOLDN,
      C => GRLFPC2_0_COMB_UN6_IUEXEC,
      Y => GRLFPC2_0_V_I_V_1_SQMUXA);
  x_grlfpc2_0_v_state_1_sqmuxa: CM8 port map (
      D0 => rst,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_V_STATE_1_SQMUXA_CM8I,
      S01 => cpi_dbg_data(28),
      S10 => NN_2,
      S11 => NN_2,
      Y => GRLFPC2_0_V_STATE_1_SQMUXA);
  x_grlfpc2_0_v_state_1_sqmuxa_1: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_X_AFQ,
      S01 => GRLFPC2_0_COMB_QNE2,
      S10 => GRLFPC2_0_R_X_SEQERR,
      S11 => NN_2,
      Y => GRLFPC2_0_V_STATE_1_SQMUXA_1);
  x_grlfpc2_0_v_state_1_sqmuxa_cm8i: CM8INV port map (
      A => GRLFPC2_0_COMB_V_FSR_TEM_1_SN_N_3,
      Y => GRLFPC2_0_V_STATE_1_SQMUXA_CM8I);
  x_grlfpc2_0_wraddr_0_sqmuxa: AND3A port map (
      A => cpi_dbg_fsr,
      B => cpi_dbg_enable,
      C => cpi_dbg_write,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA);
  x_grlfpc2_0_wraddr_0_sqmuxa_0: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_0);
  x_grlfpc2_0_wraddr_0_sqmuxa_0_0: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_0_0);
  x_grlfpc2_0_wraddr_0_sqmuxa_1: AND3B port map (
      A => GRLFPC2_0_R_X_AFSR,
      B => GRLFPC2_0_COMB_UN1_FPCI,
      C => GRLFPC2_0_R_X_LD,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_0: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_0);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_0_0: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_1: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_1);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_2: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_2);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_3: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_3);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_4: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_4);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_5: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_5);
  x_grlfpc2_0_wraddr_0_sqmuxa_1_6: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_1_6);
  x_grlfpc2_0_wraddr_0_sqmuxa_2: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_2);
  x_grlfpc2_0_wraddr_0_sqmuxa_3: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_3);
  x_grlfpc2_0_wraddr_0_sqmuxa_4: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_4);
  x_grlfpc2_0_wraddr_0_sqmuxa_5: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_5);
  x_grlfpc2_0_wraddr_0_sqmuxa_6: BUFF port map (
      A => GRLFPC2_0_WRADDR_0_SQMUXA_0_0,
      Y => GRLFPC2_0_WRADDR_0_SQMUXA_6);
  x_grlfpc2_0_wraddr_1_1x: CM8 port map (
      D0 => cpi_x_inst(26),
      D1 => cpi_dbg_addr(1),
      D2 => GRLFPC2_0_R_I_INST(26),
      D3 => cpi_dbg_addr(1),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S11 => NN_2,
      Y => RFI2_WRADDR_0_INT_13_INT_26);
  x_grlfpc2_0_wraddr_1_2x: CM8 port map (
      D0 => cpi_x_inst(27),
      D1 => cpi_dbg_addr(2),
      D2 => GRLFPC2_0_R_I_INST(27),
      D3 => cpi_dbg_addr(2),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S11 => NN_2,
      Y => RFI2_WRADDR_1_INT_14_INT_27);
  x_grlfpc2_0_wraddr_1_3x: CM8 port map (
      D0 => cpi_x_inst(28),
      D1 => cpi_dbg_addr(3),
      D2 => GRLFPC2_0_R_I_INST(28),
      D3 => cpi_dbg_addr(3),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S11 => NN_2,
      Y => RFI2_WRADDR_2_INT_15_INT_28);
  x_grlfpc2_0_wraddr_1_4x: CM8 port map (
      D0 => cpi_x_inst(29),
      D1 => cpi_dbg_addr(4),
      D2 => GRLFPC2_0_R_I_INST(29),
      D3 => cpi_dbg_addr(4),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S11 => NN_2,
      Y => RFI2_WRADDR_3_INT_16_INT_29);
  x_grlfpc2_0_wraddr_1_sqmuxa: CM8 port map (
      D0 => NN_4,
      D1 => GRLFPC2_0_R_I_EXEC,
      D2 => NN_2,
      D3 => NN_2,
      S00 => GRLFPC2_0_R_I_V,
      S01 => GRLFPC2_0_R_X_FPOP,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => GRLFPC2_0_WRADDR_1_SQMUXA);
  x_grlfpc2_0_wrdata_0x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(0),
      D1 => cpi_dbg_data(0),
      D2 => cpi_lddata(0),
      D3 => cpi_dbg_data(0),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(0));
  x_grlfpc2_0_wrdata_1x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(1),
      D1 => cpi_dbg_data(1),
      D2 => cpi_lddata(1),
      D3 => cpi_dbg_data(1),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(1));
  x_grlfpc2_0_wrdata_2x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(2),
      D1 => cpi_dbg_data(2),
      D2 => cpi_lddata(2),
      D3 => cpi_dbg_data(2),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(2));
  x_grlfpc2_0_wrdata_3x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(3),
      D1 => cpi_dbg_data(3),
      D2 => cpi_lddata(3),
      D3 => cpi_dbg_data(3),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(3));
  x_grlfpc2_0_wrdata_4x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(4),
      D1 => cpi_dbg_data(4),
      D2 => cpi_lddata(4),
      D3 => cpi_dbg_data(4),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(4));
  x_grlfpc2_0_wrdata_5x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(5),
      D1 => cpi_dbg_data(5),
      D2 => cpi_lddata(5),
      D3 => cpi_dbg_data(5),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(5));
  x_grlfpc2_0_wrdata_6x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(6),
      D1 => cpi_dbg_data(6),
      D2 => cpi_lddata(6),
      D3 => cpi_dbg_data(6),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(6));
  x_grlfpc2_0_wrdata_7x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(7),
      D1 => cpi_dbg_data(7),
      D2 => cpi_lddata(7),
      D3 => cpi_dbg_data(7),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0_0,
      S11 => NN_2,
      Y => rfi2_wrdata(7));
  x_grlfpc2_0_wrdata_8x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(8),
      D1 => cpi_dbg_data(8),
      D2 => cpi_lddata(8),
      D3 => cpi_dbg_data(8),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(8));
  x_grlfpc2_0_wrdata_9x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(9),
      D1 => cpi_dbg_data(9),
      D2 => cpi_lddata(9),
      D3 => cpi_dbg_data(9),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(9));
  x_grlfpc2_0_wrdata_10x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(10),
      D1 => cpi_dbg_data(10),
      D2 => cpi_lddata(10),
      D3 => cpi_dbg_data(10),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(10));
  x_grlfpc2_0_wrdata_11x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(11),
      D1 => cpi_dbg_data(11),
      D2 => cpi_lddata(11),
      D3 => cpi_dbg_data(11),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_1_0,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(11));
  x_grlfpc2_0_wrdata_12x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(12),
      D1 => cpi_dbg_data(12),
      D2 => cpi_lddata(12),
      D3 => cpi_dbg_data(12),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(12));
  x_grlfpc2_0_wrdata_13x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(13),
      D1 => cpi_dbg_data(13),
      D2 => cpi_lddata(13),
      D3 => cpi_dbg_data(13),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(13));
  x_grlfpc2_0_wrdata_14x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(14),
      D1 => cpi_dbg_data(14),
      D2 => cpi_lddata(14),
      D3 => cpi_dbg_data(14),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(14));
  x_grlfpc2_0_wrdata_15x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(15),
      D1 => cpi_dbg_data(15),
      D2 => cpi_lddata(15),
      D3 => cpi_dbg_data(15),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(15));
  x_grlfpc2_0_wrdata_16x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(16),
      D1 => cpi_dbg_data(16),
      D2 => cpi_lddata(16),
      D3 => cpi_dbg_data(16),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_1,
      S11 => NN_2,
      Y => rfi2_wrdata(16));
  x_grlfpc2_0_wrdata_17x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(17),
      D1 => cpi_dbg_data(17),
      D2 => cpi_lddata(17),
      D3 => cpi_dbg_data(17),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(17));
  x_grlfpc2_0_wrdata_18x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(18),
      D1 => cpi_dbg_data(18),
      D2 => cpi_lddata(18),
      D3 => cpi_dbg_data(18),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(18));
  x_grlfpc2_0_wrdata_19x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(19),
      D1 => cpi_dbg_data(19),
      D2 => cpi_lddata(19),
      D3 => cpi_dbg_data(19),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(19));
  x_grlfpc2_0_wrdata_20x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(20),
      D1 => cpi_dbg_data(20),
      D2 => cpi_lddata(20),
      D3 => cpi_dbg_data(20),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_2,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(20));
  x_grlfpc2_0_wrdata_21x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(21),
      D1 => cpi_dbg_data(21),
      D2 => cpi_lddata(21),
      D3 => cpi_dbg_data(21),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(21));
  x_grlfpc2_0_wrdata_22x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(22),
      D1 => cpi_dbg_data(22),
      D2 => cpi_lddata(22),
      D3 => cpi_dbg_data(22),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(22));
  x_grlfpc2_0_wrdata_23x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(23),
      D1 => cpi_dbg_data(23),
      D2 => cpi_lddata(23),
      D3 => cpi_dbg_data(23),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(23));
  x_grlfpc2_0_wrdata_24x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(24),
      D1 => cpi_dbg_data(24),
      D2 => cpi_lddata(24),
      D3 => cpi_dbg_data(24),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(24));
  x_grlfpc2_0_wrdata_25x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(25),
      D1 => cpi_dbg_data(25),
      D2 => cpi_lddata(25),
      D3 => cpi_dbg_data(25),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_2,
      S11 => NN_2,
      Y => rfi2_wrdata(25));
  x_grlfpc2_0_wrdata_26x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(26),
      D1 => cpi_dbg_data(26),
      D2 => cpi_lddata(26),
      D3 => cpi_dbg_data(26),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi2_wrdata(26));
  x_grlfpc2_0_wrdata_27x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(27),
      D1 => cpi_dbg_data(27),
      D2 => cpi_lddata(27),
      D3 => cpi_dbg_data(27),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi2_wrdata(27));
  x_grlfpc2_0_wrdata_28x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(28),
      D1 => cpi_dbg_data(28),
      D2 => cpi_lddata(28),
      D3 => cpi_dbg_data(28),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi2_wrdata(28));
  x_grlfpc2_0_wrdata_29x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(29),
      D1 => cpi_dbg_data(29),
      D2 => cpi_lddata(29),
      D3 => cpi_dbg_data(29),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi2_wrdata(29));
  x_grlfpc2_0_wrdata_30x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(30),
      D1 => cpi_dbg_data(30),
      D2 => cpi_lddata(30),
      D3 => cpi_dbg_data(30),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi2_wrdata(30));
  x_grlfpc2_0_wrdata_31x: CM8 port map (
      D0 => RFI1_WRDATA_31_INT_17,
      D1 => GRLFPC2_0_R_I_RES(31),
      D2 => RFI1_WRDATA_31_INT_17,
      D3 => RFI1_WRDATA_31_INT_17,
      S00 => GRLFPC2_0_COMB_RDD_3,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      Y => rfi2_wrdata(31));
  x_grlfpc2_0_wrdata_32x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(32),
      D1 => cpi_dbg_data(0),
      D2 => cpi_lddata(0),
      D3 => cpi_dbg_data(0),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi1_wrdata(0));
  x_grlfpc2_0_wrdata_33x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(33),
      D1 => cpi_dbg_data(1),
      D2 => cpi_lddata(1),
      D3 => cpi_dbg_data(1),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi1_wrdata(1));
  x_grlfpc2_0_wrdata_34x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(34),
      D1 => cpi_dbg_data(2),
      D2 => cpi_lddata(2),
      D3 => cpi_dbg_data(2),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_3,
      S11 => NN_2,
      Y => rfi1_wrdata(2));
  x_grlfpc2_0_wrdata_35x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(35),
      D1 => cpi_dbg_data(3),
      D2 => cpi_lddata(3),
      D3 => cpi_dbg_data(3),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(3));
  x_grlfpc2_0_wrdata_36x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(36),
      D1 => cpi_dbg_data(4),
      D2 => cpi_lddata(4),
      D3 => cpi_dbg_data(4),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(4));
  x_grlfpc2_0_wrdata_37x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(37),
      D1 => cpi_dbg_data(5),
      D2 => cpi_lddata(5),
      D3 => cpi_dbg_data(5),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(5));
  x_grlfpc2_0_wrdata_38x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(38),
      D1 => cpi_dbg_data(6),
      D2 => cpi_lddata(6),
      D3 => cpi_dbg_data(6),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(6));
  x_grlfpc2_0_wrdata_39x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(39),
      D1 => cpi_dbg_data(7),
      D2 => cpi_lddata(7),
      D3 => cpi_dbg_data(7),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(7));
  x_grlfpc2_0_wrdata_40x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(40),
      D1 => cpi_dbg_data(8),
      D2 => cpi_lddata(8),
      D3 => cpi_dbg_data(8),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(8));
  x_grlfpc2_0_wrdata_41x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(41),
      D1 => cpi_dbg_data(9),
      D2 => cpi_lddata(9),
      D3 => cpi_dbg_data(9),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(9));
  x_grlfpc2_0_wrdata_42x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(42),
      D1 => cpi_dbg_data(10),
      D2 => cpi_lddata(10),
      D3 => cpi_dbg_data(10),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(10));
  x_grlfpc2_0_wrdata_43x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(43),
      D1 => cpi_dbg_data(11),
      D2 => cpi_lddata(11),
      D3 => cpi_dbg_data(11),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_4,
      S11 => NN_2,
      Y => rfi1_wrdata(11));
  x_grlfpc2_0_wrdata_44x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(44),
      D1 => cpi_dbg_data(12),
      D2 => cpi_lddata(12),
      D3 => cpi_dbg_data(12),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(12));
  x_grlfpc2_0_wrdata_45x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(45),
      D1 => cpi_dbg_data(13),
      D2 => cpi_lddata(13),
      D3 => cpi_dbg_data(13),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(13));
  x_grlfpc2_0_wrdata_46x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(46),
      D1 => cpi_dbg_data(14),
      D2 => cpi_lddata(14),
      D3 => cpi_dbg_data(14),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(14));
  x_grlfpc2_0_wrdata_47x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(47),
      D1 => cpi_dbg_data(15),
      D2 => cpi_lddata(15),
      D3 => cpi_dbg_data(15),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_5,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(15));
  x_grlfpc2_0_wrdata_48x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(48),
      D1 => cpi_dbg_data(16),
      D2 => cpi_lddata(16),
      D3 => cpi_dbg_data(16),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(16));
  x_grlfpc2_0_wrdata_49x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(49),
      D1 => cpi_dbg_data(17),
      D2 => cpi_lddata(17),
      D3 => cpi_dbg_data(17),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(17));
  x_grlfpc2_0_wrdata_50x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(50),
      D1 => cpi_dbg_data(18),
      D2 => cpi_lddata(18),
      D3 => cpi_dbg_data(18),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(18));
  x_grlfpc2_0_wrdata_51x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(51),
      D1 => cpi_dbg_data(19),
      D2 => cpi_lddata(19),
      D3 => cpi_dbg_data(19),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(19));
  x_grlfpc2_0_wrdata_52x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(52),
      D1 => cpi_dbg_data(20),
      D2 => cpi_lddata(20),
      D3 => cpi_dbg_data(20),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_5,
      S11 => NN_2,
      Y => rfi1_wrdata(20));
  x_grlfpc2_0_wrdata_53x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(53),
      D1 => cpi_dbg_data(21),
      D2 => cpi_lddata(21),
      D3 => cpi_dbg_data(21),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(21));
  x_grlfpc2_0_wrdata_54x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(54),
      D1 => cpi_dbg_data(22),
      D2 => cpi_lddata(22),
      D3 => cpi_dbg_data(22),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(22));
  x_grlfpc2_0_wrdata_55x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(55),
      D1 => cpi_dbg_data(23),
      D2 => cpi_lddata(23),
      D3 => cpi_dbg_data(23),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(23));
  x_grlfpc2_0_wrdata_56x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(56),
      D1 => cpi_dbg_data(24),
      D2 => cpi_lddata(24),
      D3 => cpi_dbg_data(24),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA_6,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(24));
  x_grlfpc2_0_wrdata_57x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(57),
      D1 => cpi_dbg_data(25),
      D2 => cpi_lddata(25),
      D3 => cpi_dbg_data(25),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(25));
  x_grlfpc2_0_wrdata_58x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(58),
      D1 => cpi_dbg_data(26),
      D2 => cpi_lddata(26),
      D3 => cpi_dbg_data(26),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(26));
  x_grlfpc2_0_wrdata_59x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(59),
      D1 => cpi_dbg_data(27),
      D2 => cpi_lddata(27),
      D3 => cpi_dbg_data(27),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(27));
  x_grlfpc2_0_wrdata_60x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(60),
      D1 => cpi_dbg_data(28),
      D2 => cpi_lddata(28),
      D3 => cpi_dbg_data(28),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(28));
  x_grlfpc2_0_wrdata_61x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(61),
      D1 => cpi_dbg_data(29),
      D2 => cpi_lddata(29),
      D3 => cpi_dbg_data(29),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1_6,
      S11 => NN_2,
      Y => rfi1_wrdata(29));
  x_grlfpc2_0_wrdata_62x: CM8 port map (
      D0 => GRLFPC2_0_COMB_WRDATA_4(62),
      D1 => cpi_dbg_data(30),
      D2 => cpi_lddata(30),
      D3 => cpi_dbg_data(30),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      S11 => NN_2,
      Y => rfi1_wrdata(30));
  x_grlfpc2_0_wrdata_63x: CM8 port map (
      D0 => GRLFPC2_0_R_I_RES(63),
      D1 => cpi_dbg_data(31),
      D2 => cpi_lddata(31),
      D3 => cpi_dbg_data(31),
      S00 => GRLFPC2_0_WRADDR_0_SQMUXA,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
      S11 => NN_2,
      Y => RFI1_WRDATA_31_INT_17);
  x_grlfpc2_0_wren1_0_sqmuxa_2: AND2 port map (
      A => GRLFPC2_0_COMB_WRRES4,
      B => GRLFPC2_0_COMB_RDD_3,
      Y => GRLFPC2_0_WREN1_0_SQMUXA_2);
  x_grlfpc2_0_wren1_0_sqmuxa_3: CM8 port map (
      D0 => NN_4,
      D1 => NN_2,
      D2 => GRLFPC2_0_UN1_FPCI_3_0,
      D3 => NN_2,
      S00 => GRLFPC2_0_COMB_WRRES4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WREN2_2_SQMUXA_0,
      S11 => NN_2,
      Y => GRLFPC2_0_WREN1_0_SQMUXA_3);
  x_grlfpc2_0_wren1_m_0x: CM8 port map (
      D0 => NN_2,
      D1 => NN_2,
      D2 => GRLFPC2_0_COMB_WRRES4,
      D3 => NN_2,
      S00 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S01 => GRLFPC2_0_R_I_INST(25),
      S10 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S11 => GRLFPC2_0_WREN1_M_CM8I(0),
      Y => GRLFPC2_0_WREN1_M(0));
  x_grlfpc2_0_wren1_m_cm8i_0x: CM8INV port map (
      A => cpi_x_inst(25),
      Y => GRLFPC2_0_WREN1_M_CM8I(0));
  x_grlfpc2_0_wren1_m_n_0x: CM8 port map (
      D0 => NN_4,
      D1 => cpi_x_inst(25),
      D2 => NN_4,
      D3 => GRLFPC2_0_R_I_INST(25),
      S00 => GRLFPC2_0_COMB_WRRES4,
      S01 => NN_4,
      S10 => GRLFPC2_0_WRADDR_1_SQMUXA,
      S11 => NN_2,
      Y => GRLFPC2_0_WREN1_M_N(0));
  x_grlfpc2_0_wren2_2_sqmuxa_0: AND3B port map (
      A => GRLFPC2_0_UN1_FPCI_3_1,
      B => GRLFPC2_0_R_X_AFSR,
      C => GRLFPC2_0_R_X_LD,
      Y => GRLFPC2_0_WREN2_2_SQMUXA_0);
  x_grlfpc2_0_wren210_m_n_340x: OR3A port map (
      A => GRLFPC2_0_WREN2_2_SQMUXA_0,
      B => cpi_x_inst(25),
      C => cpi_x_inst(20),
      Y => GRLFPC2_0_WREN210_M_N(340));
  x_holdn_0: BUFF port map (
      A => holdn,
      Y => HOLDN_0);
  x_holdn_1: BUFF port map (
      A => holdn,
      Y => HOLDN_1);
  cpo_exc <= CPO_EXC_INT_1;
  cpo_cc(0) <= CPO_CC_0_INT_2;
  cpo_cc(1) <= CPO_CC_1_INT_3;
  cpo_holdn <= CPO_HOLDN_INT_4;
  rfi1_rd1addr(0) <= RFI2_RD1ADDR_0_INT_5_INT_18;
  rfi1_rd1addr(1) <= RFI2_RD1ADDR_1_INT_6_INT_19;
  rfi1_rd1addr(2) <= RFI2_RD1ADDR_2_INT_7_INT_20;
  rfi1_rd1addr(3) <= RFI2_RD1ADDR_3_INT_8_INT_21;
  rfi1_rd2addr(0) <= RFI2_RD2ADDR_0_INT_9_INT_22;
  rfi1_rd2addr(1) <= RFI2_RD2ADDR_1_INT_10_INT_23;
  rfi1_rd2addr(2) <= RFI2_RD2ADDR_2_INT_11_INT_24;
  rfi1_rd2addr(3) <= RFI2_RD2ADDR_3_INT_12_INT_25;
  rfi1_wraddr(0) <= RFI2_WRADDR_0_INT_13_INT_26;
  rfi1_wraddr(1) <= RFI2_WRADDR_1_INT_14_INT_27;
  rfi1_wraddr(2) <= RFI2_WRADDR_2_INT_15_INT_28;
  rfi1_wraddr(3) <= RFI2_WRADDR_3_INT_16_INT_29;
  rfi1_wrdata(31) <= RFI1_WRDATA_31_INT_17;
  rfi2_rd1addr(0) <= RFI2_RD1ADDR_0_INT_5_INT_18;
  rfi2_rd1addr(1) <= RFI2_RD1ADDR_1_INT_6_INT_19;
  rfi2_rd1addr(2) <= RFI2_RD1ADDR_2_INT_7_INT_20;
  rfi2_rd1addr(3) <= RFI2_RD1ADDR_3_INT_8_INT_21;
  rfi2_rd2addr(0) <= RFI2_RD2ADDR_0_INT_9_INT_22;
  rfi2_rd2addr(1) <= RFI2_RD2ADDR_1_INT_10_INT_23;
  rfi2_rd2addr(2) <= RFI2_RD2ADDR_2_INT_11_INT_24;
  rfi2_rd2addr(3) <= RFI2_RD2ADDR_3_INT_12_INT_25;
  rfi2_wraddr(0) <= RFI2_WRADDR_0_INT_13_INT_26;
  rfi2_wraddr(1) <= RFI2_WRADDR_1_INT_14_INT_27;
  rfi2_wraddr(2) <= RFI2_WRADDR_2_INT_15_INT_28;
  rfi2_wraddr(3) <= RFI2_WRADDR_3_INT_16_INT_29;
end beh;

